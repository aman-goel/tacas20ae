// RTL (Verilog) generated @ Wed Jan 31 20:28:21 2018 by V3 
//               compiled @ Jan 31 2018 12:00:50
// Internal nets are renamed with prefix "v3_1517448501_".

// Module needham
module needham
(
   v3_clock,
   f129,
   f126,
   f123,
   f119,
   f115,
   f111,
   f000,
   f130,
   f127,
   f124,
   f120,
   f116,
   f112,
   f002,
   f131,
   f128,
   f125,
   f121,
   f117,
   f113,
   f004,
   f144,
   f140,
   f136,
   f132,
   f108,
   f105,
   f102,
   f099,
   f096,
   f093,
   f090,
   f087,
   f084,
   f081,
   f078,
   f075,
   f072,
   f069,
   f066,
   f063,
   f060,
   f057,
   f054,
   f051,
   f048,
   f044,
   f040,
   f036,
   f006,
   f145,
   f141,
   f137,
   f133,
   f109,
   f106,
   f103,
   f100,
   f097,
   f094,
   f091,
   f088,
   f085,
   f082,
   f079,
   f076,
   f073,
   f070,
   f067,
   f064,
   f061,
   f058,
   f055,
   f052,
   f049,
   f045,
   f041,
   f037,
   f010,
   f146,
   f142,
   f138,
   f134,
   f110,
   f107,
   f104,
   f101,
   f098,
   f095,
   f092,
   f089,
   f086,
   f083,
   f080,
   f077,
   f074,
   f071,
   f068,
   f065,
   f062,
   f059,
   f056,
   f053,
   f050,
   f046,
   f042,
   f038,
   f014,
   f031,
   f021,
   f032,
   f022,
   f027,
   f026,
   f034,
   f024,
   f143,
   f139,
   f135,
   f122,
   f118,
   f114,
   f047,
   f043,
   f039,
   f001,
   f003,
   f005,
   f007,
   f008,
   f009,
   f011,
   f012,
   f013,
   f015,
   f016,
   f017,
   f018,
   f025,
   f028,
   f033,
   f035,
   f019,
   f020,
   f023,
   f029,
   f030,
   id78
);

   // Clock Signal for Synchronous DFF
   input v3_clock;

   // I/O Declarations
   input f129;
   input f126;
   input f123;
   input f119;
   input f115;
   input f111;
   input f000;
   input f130;
   input f127;
   input f124;
   input f120;
   input f116;
   input f112;
   input f002;
   input f131;
   input f128;
   input f125;
   input f121;
   input f117;
   input f113;
   input f004;
   input f144;
   input f140;
   input f136;
   input f132;
   input f108;
   input f105;
   input f102;
   input f099;
   input f096;
   input f093;
   input f090;
   input f087;
   input f084;
   input f081;
   input f078;
   input f075;
   input f072;
   input f069;
   input f066;
   input f063;
   input f060;
   input f057;
   input f054;
   input f051;
   input f048;
   input f044;
   input f040;
   input f036;
   input f006;
   input f145;
   input f141;
   input f137;
   input f133;
   input f109;
   input f106;
   input f103;
   input f100;
   input f097;
   input f094;
   input f091;
   input f088;
   input f085;
   input f082;
   input f079;
   input f076;
   input f073;
   input f070;
   input f067;
   input f064;
   input f061;
   input f058;
   input f055;
   input f052;
   input f049;
   input f045;
   input f041;
   input f037;
   input f010;
   input f146;
   input f142;
   input f138;
   input f134;
   input f110;
   input f107;
   input f104;
   input f101;
   input f098;
   input f095;
   input f092;
   input f089;
   input f086;
   input f083;
   input f080;
   input f077;
   input f074;
   input f071;
   input f068;
   input f065;
   input f062;
   input f059;
   input f056;
   input f053;
   input f050;
   input f046;
   input f042;
   input f038;
   input f014;
   input f031;
   input f021;
   input f032;
   input f022;
   input f027;
   input f026;
   input f034;
   input f024;
   input f143;
   input f139;
   input f135;
   input f122;
   input f118;
   input f114;
   input f047;
   input f043;
   input f039;
   input f001;
   input f003;
   input f005;
   input f007;
   input f008;
   input f009;
   input f011;
   input f012;
   input f013;
   input f015;
   input f016;
   input f017;
   input f018;
   input f025;
   input f028;
   input f033;
   input f035;
   input f019;
   input f020;
   input f023;
   input f029;
   input f030;
   output id78;

   // Wire and Reg Declarations
   wire id0;
   reg [15:0] v_m_initiator_0 = 0;
   reg [15:0] v_party_nonce_initiator_0 = 0;
   reg [15:0] v_m_initiator_1 = 0;
   reg [15:0] v_party_nonce_initiator_1 = 0;
   reg [15:0] v_m_initiator_2 = 0;
   reg [15:0] v_party_nonce_initiator_2 = 0;
   reg [15:0] v_m_responder_0 = 0;
   reg [15:0] v_party_responder_0 = 0;
   reg [15:0] v_party_nonce_responder_0 = 0;
   reg [15:0] v_m_responder_1 = 0;
   reg [15:0] v_party_responder_1 = 0;
   reg [15:0] v_party_nonce_responder_1 = 0;
   reg [15:0] v_m_responder_2 = 0;
   reg [15:0] v_party_responder_2 = 0;
   reg [15:0] v_party_nonce_responder_2 = 0;
   reg [7:0] v_kNa = 0;
   reg [7:0] v_kNb = 0;
   reg [7:0] v_k_Na_Nb__A = 0;
   reg [7:0] v_k_Na_A__B = 0;
   reg [7:0] v_k_Nb__B = 0;
   reg [15:0] v_m_intruder = 0;
   reg a_start_initiator_0 = 0;
   reg a_wait_resp_initiator_0 = 0;
   reg a_got_resp_initiator_0 = 0;
   reg a_commited_initiator_0 = 0;
   reg a_finished_initiator_0 = 0;
   reg a_corrupted_initiator_0 = 0;
   reg a_start_initiator_1 = 0;
   reg a_wait_resp_initiator_1 = 0;
   reg a_got_resp_initiator_1 = 0;
   reg a_commited_initiator_1 = 0;
   reg a_finished_initiator_1 = 0;
   reg a_corrupted_initiator_1 = 0;
   reg a_start_initiator_2 = 0;
   reg a_wait_resp_initiator_2 = 0;
   reg a_got_resp_initiator_2 = 0;
   reg a_commited_initiator_2 = 0;
   reg a_finished_initiator_2 = 0;
   reg a_corrupted_initiator_2 = 0;
   reg a_start_responder_0 = 0;
   reg a_got_msg_responder_0 = 0;
   reg a_send_reply_responder_0 = 0;
   reg a_wait_resp_responder_0 = 0;
   reg a_got_resp_responder_0 = 0;
   reg a_finished_responder_0 = 0;
   reg a_corrupted_responder_0 = 0;
   reg a_start_responder_1 = 0;
   reg a_got_msg_responder_1 = 0;
   reg a_send_reply_responder_1 = 0;
   reg a_wait_resp_responder_1 = 0;
   reg a_got_resp_responder_1 = 0;
   reg a_finished_responder_1 = 0;
   reg a_corrupted_responder_1 = 0;
   reg a_start_responder_2 = 0;
   reg a_got_msg_responder_2 = 0;
   reg a_send_reply_responder_2 = 0;
   reg a_wait_resp_responder_2 = 0;
   reg a_got_resp_responder_2 = 0;
   reg a_finished_responder_2 = 0;
   reg a_corrupted_responder_2 = 0;
   reg a_q = 0;
   reg a_got3 = 0;
   reg a_c1 = 0;
   reg a_c2 = 0;
   reg a_d1 = 0;
   reg a_got2 = 0;
   reg a_e1 = 0;
   reg a_f1 = 0;
   reg dve_invalid = 0;
   wire [31:0] v3_1517448501_70;
   wire [15:0] v3_1517448501_71;
   wire [31:0] v3_1517448501_72;
   wire [4:0] v3_1517448501_73;
   wire [31:0] v3_1517448501_74;
   wire [31:0] v3_1517448501_75;
   wire [31:0] v3_1517448501_76;
   wire v3_1517448501_77;
   wire v3_1517448501_78;
   wire v3_1517448501_79;
   wire v3_1517448501_80;
   wire f129;
   wire [15:0] v3_1517448501_82;
   wire f126;
   wire [15:0] v3_1517448501_84;
   wire f123;
   wire [15:0] v3_1517448501_86;
   wire f119;
   wire [31:0] v3_1517448501_88;
   wire [31:0] v3_1517448501_89;
   wire [31:0] v3_1517448501_90;
   wire [31:0] v3_1517448501_91;
   wire [31:0] v3_1517448501_92;
   wire v3_1517448501_93;
   wire [31:0] v3_1517448501_94;
   wire [31:0] v3_1517448501_95;
   wire [31:0] v3_1517448501_96;
   wire [31:0] v3_1517448501_97;
   wire [31:0] v3_1517448501_98;
   wire [31:0] v3_1517448501_99;
   wire v3_1517448501_100;
   wire [31:0] v3_1517448501_101;
   wire [31:0] v3_1517448501_102;
   wire [31:0] v3_1517448501_103;
   wire [15:0] v3_1517448501_104;
   wire f115;
   wire [31:0] v3_1517448501_106;
   wire [31:0] v3_1517448501_107;
   wire [31:0] v3_1517448501_108;
   wire [31:0] v3_1517448501_109;
   wire [31:0] v3_1517448501_110;
   wire v3_1517448501_111;
   wire [31:0] v3_1517448501_112;
   wire [31:0] v3_1517448501_113;
   wire [31:0] v3_1517448501_114;
   wire [31:0] v3_1517448501_115;
   wire [31:0] v3_1517448501_116;
   wire v3_1517448501_117;
   wire [31:0] v3_1517448501_118;
   wire [31:0] v3_1517448501_119;
   wire [31:0] v3_1517448501_120;
   wire [15:0] v3_1517448501_121;
   wire f111;
   wire [31:0] v3_1517448501_123;
   wire [31:0] v3_1517448501_124;
   wire [31:0] v3_1517448501_125;
   wire [31:0] v3_1517448501_126;
   wire [31:0] v3_1517448501_127;
   wire v3_1517448501_128;
   wire [31:0] v3_1517448501_129;
   wire [31:0] v3_1517448501_130;
   wire [31:0] v3_1517448501_131;
   wire [31:0] v3_1517448501_132;
   wire [15:0] v3_1517448501_133;
   wire [15:0] v3_1517448501_134;
   wire [15:0] v3_1517448501_135;
   wire [15:0] v3_1517448501_136;
   wire [15:0] v3_1517448501_137;
   wire [15:0] v3_1517448501_138;
   wire [15:0] v3_1517448501_139;
   wire [15:0] v3_1517448501_140;
   wire f000;
   wire [31:0] v3_1517448501_142;
   wire [31:0] v3_1517448501_143;
   wire [31:0] v3_1517448501_144;
   wire [31:0] v3_1517448501_145;
   wire v3_1517448501_146;
   wire [31:0] v3_1517448501_147;
   wire [31:0] v3_1517448501_148;
   wire v3_1517448501_149;
   wire v3_1517448501_150;
   wire [31:0] v3_1517448501_151;
   wire [31:0] v3_1517448501_152;
   wire [31:0] v3_1517448501_153;
   wire [31:0] v3_1517448501_154;
   wire [31:0] v3_1517448501_155;
   wire [31:0] v3_1517448501_156;
   wire [31:0] v3_1517448501_157;
   wire [31:0] v3_1517448501_158;
   wire v3_1517448501_159;
   wire v3_1517448501_160;
   wire v3_1517448501_161;
   wire [31:0] v3_1517448501_162;
   wire [31:0] v3_1517448501_163;
   wire [31:0] v3_1517448501_164;
   wire [31:0] v3_1517448501_165;
   wire [31:0] v3_1517448501_166;
   wire [31:0] v3_1517448501_167;
   wire [31:0] v3_1517448501_168;
   wire [15:0] v3_1517448501_169;
   wire [15:0] v3_1517448501_170;
   wire [15:0] v3_1517448501_171;
   wire f130;
   wire f127;
   wire f124;
   wire f120;
   wire f116;
   wire f112;
   wire [15:0] v3_1517448501_178;
   wire [15:0] v3_1517448501_179;
   wire [15:0] v3_1517448501_180;
   wire [15:0] v3_1517448501_181;
   wire [15:0] v3_1517448501_182;
   wire [15:0] v3_1517448501_183;
   wire [15:0] v3_1517448501_184;
   wire f002;
   wire [31:0] v3_1517448501_186;
   wire [31:0] v3_1517448501_187;
   wire [31:0] v3_1517448501_188;
   wire [31:0] v3_1517448501_189;
   wire v3_1517448501_190;
   wire [31:0] v3_1517448501_191;
   wire v3_1517448501_192;
   wire v3_1517448501_193;
   wire [31:0] v3_1517448501_194;
   wire [31:0] v3_1517448501_195;
   wire [31:0] v3_1517448501_196;
   wire [31:0] v3_1517448501_197;
   wire [31:0] v3_1517448501_198;
   wire [31:0] v3_1517448501_199;
   wire [31:0] v3_1517448501_200;
   wire [31:0] v3_1517448501_201;
   wire v3_1517448501_202;
   wire v3_1517448501_203;
   wire v3_1517448501_204;
   wire [31:0] v3_1517448501_205;
   wire [31:0] v3_1517448501_206;
   wire [31:0] v3_1517448501_207;
   wire [31:0] v3_1517448501_208;
   wire [31:0] v3_1517448501_209;
   wire [31:0] v3_1517448501_210;
   wire [31:0] v3_1517448501_211;
   wire [15:0] v3_1517448501_212;
   wire [15:0] v3_1517448501_213;
   wire [15:0] v3_1517448501_214;
   wire f131;
   wire f128;
   wire f125;
   wire f121;
   wire f117;
   wire f113;
   wire [15:0] v3_1517448501_221;
   wire [15:0] v3_1517448501_222;
   wire [15:0] v3_1517448501_223;
   wire [15:0] v3_1517448501_224;
   wire [15:0] v3_1517448501_225;
   wire [15:0] v3_1517448501_226;
   wire [15:0] v3_1517448501_227;
   wire f004;
   wire [31:0] v3_1517448501_229;
   wire [31:0] v3_1517448501_230;
   wire [31:0] v3_1517448501_231;
   wire [31:0] v3_1517448501_232;
   wire v3_1517448501_233;
   wire [31:0] v3_1517448501_234;
   wire v3_1517448501_235;
   wire v3_1517448501_236;
   wire [31:0] v3_1517448501_237;
   wire [31:0] v3_1517448501_238;
   wire [31:0] v3_1517448501_239;
   wire [31:0] v3_1517448501_240;
   wire [31:0] v3_1517448501_241;
   wire [31:0] v3_1517448501_242;
   wire [31:0] v3_1517448501_243;
   wire [31:0] v3_1517448501_244;
   wire v3_1517448501_245;
   wire v3_1517448501_246;
   wire v3_1517448501_247;
   wire [31:0] v3_1517448501_248;
   wire [31:0] v3_1517448501_249;
   wire [31:0] v3_1517448501_250;
   wire [31:0] v3_1517448501_251;
   wire [31:0] v3_1517448501_252;
   wire [31:0] v3_1517448501_253;
   wire [31:0] v3_1517448501_254;
   wire [15:0] v3_1517448501_255;
   wire [15:0] v3_1517448501_256;
   wire [15:0] v3_1517448501_257;
   wire f144;
   wire [15:0] v3_1517448501_259;
   wire f140;
   wire [31:0] v3_1517448501_261;
   wire [31:0] v3_1517448501_262;
   wire [31:0] v3_1517448501_263;
   wire [31:0] v3_1517448501_264;
   wire [31:0] v3_1517448501_265;
   wire v3_1517448501_266;
   wire [31:0] v3_1517448501_267;
   wire [15:0] v3_1517448501_268;
   wire f136;
   wire [31:0] v3_1517448501_270;
   wire [31:0] v3_1517448501_271;
   wire [31:0] v3_1517448501_272;
   wire [31:0] v3_1517448501_273;
   wire [31:0] v3_1517448501_274;
   wire v3_1517448501_275;
   wire [31:0] v3_1517448501_276;
   wire [15:0] v3_1517448501_277;
   wire f132;
   wire [31:0] v3_1517448501_279;
   wire [31:0] v3_1517448501_280;
   wire [31:0] v3_1517448501_281;
   wire [31:0] v3_1517448501_282;
   wire [31:0] v3_1517448501_283;
   wire v3_1517448501_284;
   wire [31:0] v3_1517448501_285;
   wire [15:0] v3_1517448501_286;
   wire f108;
   wire [15:0] v3_1517448501_288;
   wire f105;
   wire [15:0] v3_1517448501_290;
   wire f102;
   wire [15:0] v3_1517448501_292;
   wire f099;
   wire [15:0] v3_1517448501_294;
   wire f096;
   wire [15:0] v3_1517448501_296;
   wire f093;
   wire [15:0] v3_1517448501_298;
   wire f090;
   wire [15:0] v3_1517448501_300;
   wire f087;
   wire [15:0] v3_1517448501_302;
   wire f084;
   wire [15:0] v3_1517448501_304;
   wire f081;
   wire [15:0] v3_1517448501_306;
   wire f078;
   wire [15:0] v3_1517448501_308;
   wire f075;
   wire [15:0] v3_1517448501_310;
   wire f072;
   wire [15:0] v3_1517448501_312;
   wire f069;
   wire [15:0] v3_1517448501_314;
   wire f066;
   wire [15:0] v3_1517448501_316;
   wire f063;
   wire [15:0] v3_1517448501_318;
   wire f060;
   wire [15:0] v3_1517448501_320;
   wire f057;
   wire [15:0] v3_1517448501_322;
   wire f054;
   wire [15:0] v3_1517448501_324;
   wire f051;
   wire [15:0] v3_1517448501_326;
   wire f048;
   wire [15:0] v3_1517448501_328;
   wire f044;
   wire [15:0] v3_1517448501_330;
   wire f040;
   wire [15:0] v3_1517448501_332;
   wire f036;
   wire [15:0] v3_1517448501_334;
   wire [15:0] v3_1517448501_335;
   wire [15:0] v3_1517448501_336;
   wire [15:0] v3_1517448501_337;
   wire [15:0] v3_1517448501_338;
   wire [15:0] v3_1517448501_339;
   wire [15:0] v3_1517448501_340;
   wire [15:0] v3_1517448501_341;
   wire [15:0] v3_1517448501_342;
   wire [15:0] v3_1517448501_343;
   wire [15:0] v3_1517448501_344;
   wire [15:0] v3_1517448501_345;
   wire [15:0] v3_1517448501_346;
   wire [15:0] v3_1517448501_347;
   wire [15:0] v3_1517448501_348;
   wire [15:0] v3_1517448501_349;
   wire [15:0] v3_1517448501_350;
   wire [15:0] v3_1517448501_351;
   wire [15:0] v3_1517448501_352;
   wire [15:0] v3_1517448501_353;
   wire [15:0] v3_1517448501_354;
   wire [15:0] v3_1517448501_355;
   wire [15:0] v3_1517448501_356;
   wire [15:0] v3_1517448501_357;
   wire [15:0] v3_1517448501_358;
   wire [15:0] v3_1517448501_359;
   wire [15:0] v3_1517448501_360;
   wire [15:0] v3_1517448501_361;
   wire [15:0] v3_1517448501_362;
   wire f006;
   wire [31:0] v3_1517448501_364;
   wire [31:0] v3_1517448501_365;
   wire [31:0] v3_1517448501_366;
   wire [31:0] v3_1517448501_367;
   wire v3_1517448501_368;
   wire [31:0] v3_1517448501_369;
   wire v3_1517448501_370;
   wire v3_1517448501_371;
   wire [31:0] v3_1517448501_372;
   wire [31:0] v3_1517448501_373;
   wire [31:0] v3_1517448501_374;
   wire [31:0] v3_1517448501_375;
   wire [31:0] v3_1517448501_376;
   wire [31:0] v3_1517448501_377;
   wire [31:0] v3_1517448501_378;
   wire [31:0] v3_1517448501_379;
   wire v3_1517448501_380;
   wire v3_1517448501_381;
   wire v3_1517448501_382;
   wire [31:0] v3_1517448501_383;
   wire [31:0] v3_1517448501_384;
   wire [31:0] v3_1517448501_385;
   wire [31:0] v3_1517448501_386;
   wire [31:0] v3_1517448501_387;
   wire [31:0] v3_1517448501_388;
   wire [31:0] v3_1517448501_389;
   wire [15:0] v3_1517448501_390;
   wire [15:0] v3_1517448501_391;
   wire [15:0] v3_1517448501_392;
   wire [31:0] v3_1517448501_393;
   wire v3_1517448501_394;
   wire v3_1517448501_395;
   wire [31:0] v3_1517448501_396;
   wire [31:0] v3_1517448501_397;
   wire [31:0] v3_1517448501_398;
   wire [31:0] v3_1517448501_399;
   wire [31:0] v3_1517448501_400;
   wire [31:0] v3_1517448501_401;
   wire [31:0] v3_1517448501_402;
   wire [15:0] v3_1517448501_403;
   wire [15:0] v3_1517448501_404;
   wire [15:0] v3_1517448501_405;
   wire f145;
   wire f141;
   wire f137;
   wire f133;
   wire f109;
   wire f106;
   wire f103;
   wire f100;
   wire f097;
   wire f094;
   wire f091;
   wire f088;
   wire f085;
   wire f082;
   wire f079;
   wire f076;
   wire f073;
   wire f070;
   wire f067;
   wire f064;
   wire f061;
   wire f058;
   wire f055;
   wire f052;
   wire f049;
   wire f045;
   wire f041;
   wire f037;
   wire [15:0] v3_1517448501_434;
   wire [15:0] v3_1517448501_435;
   wire [15:0] v3_1517448501_436;
   wire [15:0] v3_1517448501_437;
   wire [15:0] v3_1517448501_438;
   wire [15:0] v3_1517448501_439;
   wire [15:0] v3_1517448501_440;
   wire [15:0] v3_1517448501_441;
   wire [15:0] v3_1517448501_442;
   wire [15:0] v3_1517448501_443;
   wire [15:0] v3_1517448501_444;
   wire [15:0] v3_1517448501_445;
   wire [15:0] v3_1517448501_446;
   wire [15:0] v3_1517448501_447;
   wire [15:0] v3_1517448501_448;
   wire [15:0] v3_1517448501_449;
   wire [15:0] v3_1517448501_450;
   wire [15:0] v3_1517448501_451;
   wire [15:0] v3_1517448501_452;
   wire [15:0] v3_1517448501_453;
   wire [15:0] v3_1517448501_454;
   wire [15:0] v3_1517448501_455;
   wire [15:0] v3_1517448501_456;
   wire [15:0] v3_1517448501_457;
   wire [15:0] v3_1517448501_458;
   wire [15:0] v3_1517448501_459;
   wire [15:0] v3_1517448501_460;
   wire [15:0] v3_1517448501_461;
   wire [15:0] v3_1517448501_462;
   wire f010;
   wire [31:0] v3_1517448501_464;
   wire [31:0] v3_1517448501_465;
   wire [31:0] v3_1517448501_466;
   wire [31:0] v3_1517448501_467;
   wire v3_1517448501_468;
   wire [31:0] v3_1517448501_469;
   wire v3_1517448501_470;
   wire v3_1517448501_471;
   wire [31:0] v3_1517448501_472;
   wire [31:0] v3_1517448501_473;
   wire [31:0] v3_1517448501_474;
   wire [31:0] v3_1517448501_475;
   wire [31:0] v3_1517448501_476;
   wire [31:0] v3_1517448501_477;
   wire [31:0] v3_1517448501_478;
   wire [31:0] v3_1517448501_479;
   wire v3_1517448501_480;
   wire v3_1517448501_481;
   wire v3_1517448501_482;
   wire [31:0] v3_1517448501_483;
   wire [31:0] v3_1517448501_484;
   wire [31:0] v3_1517448501_485;
   wire [31:0] v3_1517448501_486;
   wire [31:0] v3_1517448501_487;
   wire [31:0] v3_1517448501_488;
   wire [31:0] v3_1517448501_489;
   wire [15:0] v3_1517448501_490;
   wire [15:0] v3_1517448501_491;
   wire [15:0] v3_1517448501_492;
   wire [31:0] v3_1517448501_493;
   wire v3_1517448501_494;
   wire v3_1517448501_495;
   wire [31:0] v3_1517448501_496;
   wire [31:0] v3_1517448501_497;
   wire [31:0] v3_1517448501_498;
   wire [31:0] v3_1517448501_499;
   wire [31:0] v3_1517448501_500;
   wire [31:0] v3_1517448501_501;
   wire [31:0] v3_1517448501_502;
   wire [15:0] v3_1517448501_503;
   wire [15:0] v3_1517448501_504;
   wire [15:0] v3_1517448501_505;
   wire f146;
   wire f142;
   wire f138;
   wire f134;
   wire f110;
   wire f107;
   wire f104;
   wire f101;
   wire f098;
   wire f095;
   wire f092;
   wire f089;
   wire f086;
   wire f083;
   wire f080;
   wire f077;
   wire f074;
   wire f071;
   wire f068;
   wire f065;
   wire f062;
   wire f059;
   wire f056;
   wire f053;
   wire f050;
   wire f046;
   wire f042;
   wire f038;
   wire [15:0] v3_1517448501_534;
   wire [15:0] v3_1517448501_535;
   wire [15:0] v3_1517448501_536;
   wire [15:0] v3_1517448501_537;
   wire [15:0] v3_1517448501_538;
   wire [15:0] v3_1517448501_539;
   wire [15:0] v3_1517448501_540;
   wire [15:0] v3_1517448501_541;
   wire [15:0] v3_1517448501_542;
   wire [15:0] v3_1517448501_543;
   wire [15:0] v3_1517448501_544;
   wire [15:0] v3_1517448501_545;
   wire [15:0] v3_1517448501_546;
   wire [15:0] v3_1517448501_547;
   wire [15:0] v3_1517448501_548;
   wire [15:0] v3_1517448501_549;
   wire [15:0] v3_1517448501_550;
   wire [15:0] v3_1517448501_551;
   wire [15:0] v3_1517448501_552;
   wire [15:0] v3_1517448501_553;
   wire [15:0] v3_1517448501_554;
   wire [15:0] v3_1517448501_555;
   wire [15:0] v3_1517448501_556;
   wire [15:0] v3_1517448501_557;
   wire [15:0] v3_1517448501_558;
   wire [15:0] v3_1517448501_559;
   wire [15:0] v3_1517448501_560;
   wire [15:0] v3_1517448501_561;
   wire [15:0] v3_1517448501_562;
   wire f014;
   wire [31:0] v3_1517448501_564;
   wire [31:0] v3_1517448501_565;
   wire [31:0] v3_1517448501_566;
   wire [31:0] v3_1517448501_567;
   wire v3_1517448501_568;
   wire [31:0] v3_1517448501_569;
   wire v3_1517448501_570;
   wire v3_1517448501_571;
   wire [31:0] v3_1517448501_572;
   wire [31:0] v3_1517448501_573;
   wire [31:0] v3_1517448501_574;
   wire [31:0] v3_1517448501_575;
   wire [31:0] v3_1517448501_576;
   wire [31:0] v3_1517448501_577;
   wire [31:0] v3_1517448501_578;
   wire [31:0] v3_1517448501_579;
   wire v3_1517448501_580;
   wire v3_1517448501_581;
   wire v3_1517448501_582;
   wire [31:0] v3_1517448501_583;
   wire [31:0] v3_1517448501_584;
   wire [31:0] v3_1517448501_585;
   wire [31:0] v3_1517448501_586;
   wire [31:0] v3_1517448501_587;
   wire [31:0] v3_1517448501_588;
   wire [31:0] v3_1517448501_589;
   wire [15:0] v3_1517448501_590;
   wire [15:0] v3_1517448501_591;
   wire [15:0] v3_1517448501_592;
   wire [31:0] v3_1517448501_593;
   wire v3_1517448501_594;
   wire v3_1517448501_595;
   wire [31:0] v3_1517448501_596;
   wire [31:0] v3_1517448501_597;
   wire [31:0] v3_1517448501_598;
   wire [31:0] v3_1517448501_599;
   wire [31:0] v3_1517448501_600;
   wire [31:0] v3_1517448501_601;
   wire [31:0] v3_1517448501_602;
   wire [15:0] v3_1517448501_603;
   wire [15:0] v3_1517448501_604;
   wire [15:0] v3_1517448501_605;
   wire f031;
   wire [7:0] v3_1517448501_607;
   wire f021;
   wire [7:0] v3_1517448501_609;
   wire [7:0] v3_1517448501_610;
   wire [7:0] v3_1517448501_611;
   wire f032;
   wire f022;
   wire [7:0] v3_1517448501_614;
   wire [7:0] v3_1517448501_615;
   wire [7:0] v3_1517448501_616;
   wire f027;
   wire [7:0] v3_1517448501_618;
   wire [7:0] v3_1517448501_619;
   wire f026;
   wire [7:0] v3_1517448501_621;
   wire [7:0] v3_1517448501_622;
   wire f034;
   wire f024;
   wire [7:0] v3_1517448501_625;
   wire [7:0] v3_1517448501_626;
   wire [7:0] v3_1517448501_627;
   wire f143;
   wire f139;
   wire f135;
   wire f122;
   wire f118;
   wire f114;
   wire f047;
   wire f043;
   wire f039;
   wire [15:0] v3_1517448501_637;
   wire [15:0] v3_1517448501_638;
   wire [15:0] v3_1517448501_639;
   wire [15:0] v3_1517448501_640;
   wire [15:0] v3_1517448501_641;
   wire [15:0] v3_1517448501_642;
   wire [15:0] v3_1517448501_643;
   wire [15:0] v3_1517448501_644;
   wire [15:0] v3_1517448501_645;
   wire [15:0] v3_1517448501_646;
   wire v3_1517448501_647;
   wire v3_1517448501_648;
   wire v3_1517448501_649;
   wire v3_1517448501_650;
   wire v3_1517448501_651;
   wire v3_1517448501_652;
   wire v3_1517448501_653;
   wire v3_1517448501_654;
   wire v3_1517448501_655;
   wire v3_1517448501_656;
   wire v3_1517448501_657;
   wire v3_1517448501_658;
   wire v3_1517448501_659;
   wire v3_1517448501_660;
   wire v3_1517448501_661;
   wire v3_1517448501_662;
   wire v3_1517448501_663;
   wire v3_1517448501_664;
   wire v3_1517448501_665;
   wire v3_1517448501_666;
   wire v3_1517448501_667;
   wire f001;
   wire v3_1517448501_669;
   wire v3_1517448501_670;
   wire v3_1517448501_671;
   wire v3_1517448501_672;
   wire v3_1517448501_673;
   wire v3_1517448501_674;
   wire v3_1517448501_675;
   wire v3_1517448501_676;
   wire v3_1517448501_677;
   wire v3_1517448501_678;
   wire v3_1517448501_679;
   wire v3_1517448501_680;
   wire v3_1517448501_681;
   wire v3_1517448501_682;
   wire v3_1517448501_683;
   wire v3_1517448501_684;
   wire v3_1517448501_685;
   wire v3_1517448501_686;
   wire v3_1517448501_687;
   wire v3_1517448501_688;
   wire v3_1517448501_689;
   wire v3_1517448501_690;
   wire v3_1517448501_691;
   wire v3_1517448501_692;
   wire v3_1517448501_693;
   wire v3_1517448501_694;
   wire v3_1517448501_695;
   wire v3_1517448501_696;
   wire v3_1517448501_697;
   wire v3_1517448501_698;
   wire v3_1517448501_699;
   wire v3_1517448501_700;
   wire v3_1517448501_701;
   wire v3_1517448501_702;
   wire v3_1517448501_703;
   wire v3_1517448501_704;
   wire v3_1517448501_705;
   wire v3_1517448501_706;
   wire v3_1517448501_707;
   wire v3_1517448501_708;
   wire v3_1517448501_709;
   wire v3_1517448501_710;
   wire v3_1517448501_711;
   wire v3_1517448501_712;
   wire v3_1517448501_713;
   wire v3_1517448501_714;
   wire v3_1517448501_715;
   wire v3_1517448501_716;
   wire v3_1517448501_717;
   wire v3_1517448501_718;
   wire v3_1517448501_719;
   wire v3_1517448501_720;
   wire v3_1517448501_721;
   wire v3_1517448501_722;
   wire f003;
   wire v3_1517448501_724;
   wire v3_1517448501_725;
   wire v3_1517448501_726;
   wire v3_1517448501_727;
   wire v3_1517448501_728;
   wire v3_1517448501_729;
   wire v3_1517448501_730;
   wire v3_1517448501_731;
   wire v3_1517448501_732;
   wire v3_1517448501_733;
   wire v3_1517448501_734;
   wire v3_1517448501_735;
   wire v3_1517448501_736;
   wire v3_1517448501_737;
   wire v3_1517448501_738;
   wire v3_1517448501_739;
   wire v3_1517448501_740;
   wire v3_1517448501_741;
   wire v3_1517448501_742;
   wire v3_1517448501_743;
   wire v3_1517448501_744;
   wire v3_1517448501_745;
   wire v3_1517448501_746;
   wire v3_1517448501_747;
   wire v3_1517448501_748;
   wire v3_1517448501_749;
   wire v3_1517448501_750;
   wire v3_1517448501_751;
   wire v3_1517448501_752;
   wire v3_1517448501_753;
   wire v3_1517448501_754;
   wire v3_1517448501_755;
   wire v3_1517448501_756;
   wire v3_1517448501_757;
   wire v3_1517448501_758;
   wire v3_1517448501_759;
   wire v3_1517448501_760;
   wire v3_1517448501_761;
   wire v3_1517448501_762;
   wire v3_1517448501_763;
   wire v3_1517448501_764;
   wire v3_1517448501_765;
   wire v3_1517448501_766;
   wire v3_1517448501_767;
   wire v3_1517448501_768;
   wire v3_1517448501_769;
   wire v3_1517448501_770;
   wire v3_1517448501_771;
   wire v3_1517448501_772;
   wire v3_1517448501_773;
   wire v3_1517448501_774;
   wire v3_1517448501_775;
   wire v3_1517448501_776;
   wire v3_1517448501_777;
   wire f005;
   wire v3_1517448501_779;
   wire v3_1517448501_780;
   wire v3_1517448501_781;
   wire v3_1517448501_782;
   wire v3_1517448501_783;
   wire v3_1517448501_784;
   wire v3_1517448501_785;
   wire v3_1517448501_786;
   wire v3_1517448501_787;
   wire v3_1517448501_788;
   wire v3_1517448501_789;
   wire v3_1517448501_790;
   wire v3_1517448501_791;
   wire v3_1517448501_792;
   wire v3_1517448501_793;
   wire v3_1517448501_794;
   wire v3_1517448501_795;
   wire v3_1517448501_796;
   wire v3_1517448501_797;
   wire v3_1517448501_798;
   wire v3_1517448501_799;
   wire v3_1517448501_800;
   wire v3_1517448501_801;
   wire v3_1517448501_802;
   wire v3_1517448501_803;
   wire v3_1517448501_804;
   wire v3_1517448501_805;
   wire v3_1517448501_806;
   wire v3_1517448501_807;
   wire v3_1517448501_808;
   wire v3_1517448501_809;
   wire v3_1517448501_810;
   wire v3_1517448501_811;
   wire v3_1517448501_812;
   wire v3_1517448501_813;
   wire v3_1517448501_814;
   wire v3_1517448501_815;
   wire v3_1517448501_816;
   wire v3_1517448501_817;
   wire v3_1517448501_818;
   wire v3_1517448501_819;
   wire v3_1517448501_820;
   wire v3_1517448501_821;
   wire v3_1517448501_822;
   wire v3_1517448501_823;
   wire v3_1517448501_824;
   wire v3_1517448501_825;
   wire v3_1517448501_826;
   wire v3_1517448501_827;
   wire v3_1517448501_828;
   wire v3_1517448501_829;
   wire v3_1517448501_830;
   wire v3_1517448501_831;
   wire v3_1517448501_832;
   wire v3_1517448501_833;
   wire v3_1517448501_834;
   wire v3_1517448501_835;
   wire v3_1517448501_836;
   wire v3_1517448501_837;
   wire f007;
   wire v3_1517448501_839;
   wire v3_1517448501_840;
   wire v3_1517448501_841;
   wire v3_1517448501_842;
   wire v3_1517448501_843;
   wire v3_1517448501_844;
   wire v3_1517448501_845;
   wire v3_1517448501_846;
   wire v3_1517448501_847;
   wire v3_1517448501_848;
   wire v3_1517448501_849;
   wire v3_1517448501_850;
   wire v3_1517448501_851;
   wire v3_1517448501_852;
   wire v3_1517448501_853;
   wire v3_1517448501_854;
   wire v3_1517448501_855;
   wire v3_1517448501_856;
   wire v3_1517448501_857;
   wire v3_1517448501_858;
   wire v3_1517448501_859;
   wire v3_1517448501_860;
   wire v3_1517448501_861;
   wire v3_1517448501_862;
   wire v3_1517448501_863;
   wire v3_1517448501_864;
   wire v3_1517448501_865;
   wire v3_1517448501_866;
   wire v3_1517448501_867;
   wire v3_1517448501_868;
   wire v3_1517448501_869;
   wire v3_1517448501_870;
   wire v3_1517448501_871;
   wire v3_1517448501_872;
   wire v3_1517448501_873;
   wire v3_1517448501_874;
   wire v3_1517448501_875;
   wire v3_1517448501_876;
   wire v3_1517448501_877;
   wire v3_1517448501_878;
   wire v3_1517448501_879;
   wire v3_1517448501_880;
   wire v3_1517448501_881;
   wire v3_1517448501_882;
   wire v3_1517448501_883;
   wire v3_1517448501_884;
   wire v3_1517448501_885;
   wire v3_1517448501_886;
   wire v3_1517448501_887;
   wire v3_1517448501_888;
   wire v3_1517448501_889;
   wire v3_1517448501_890;
   wire v3_1517448501_891;
   wire v3_1517448501_892;
   wire v3_1517448501_893;
   wire v3_1517448501_894;
   wire v3_1517448501_895;
   wire v3_1517448501_896;
   wire v3_1517448501_897;
   wire v3_1517448501_898;
   wire v3_1517448501_899;
   wire v3_1517448501_900;
   wire v3_1517448501_901;
   wire v3_1517448501_902;
   wire v3_1517448501_903;
   wire v3_1517448501_904;
   wire v3_1517448501_905;
   wire v3_1517448501_906;
   wire v3_1517448501_907;
   wire v3_1517448501_908;
   wire f008;
   wire v3_1517448501_910;
   wire f009;
   wire v3_1517448501_912;
   wire v3_1517448501_913;
   wire v3_1517448501_914;
   wire v3_1517448501_915;
   wire v3_1517448501_916;
   wire v3_1517448501_917;
   wire v3_1517448501_918;
   wire v3_1517448501_919;
   wire v3_1517448501_920;
   wire v3_1517448501_921;
   wire v3_1517448501_922;
   wire v3_1517448501_923;
   wire v3_1517448501_924;
   wire v3_1517448501_925;
   wire v3_1517448501_926;
   wire v3_1517448501_927;
   wire v3_1517448501_928;
   wire v3_1517448501_929;
   wire v3_1517448501_930;
   wire v3_1517448501_931;
   wire v3_1517448501_932;
   wire v3_1517448501_933;
   wire v3_1517448501_934;
   wire v3_1517448501_935;
   wire v3_1517448501_936;
   wire v3_1517448501_937;
   wire v3_1517448501_938;
   wire v3_1517448501_939;
   wire v3_1517448501_940;
   wire v3_1517448501_941;
   wire v3_1517448501_942;
   wire v3_1517448501_943;
   wire v3_1517448501_944;
   wire v3_1517448501_945;
   wire v3_1517448501_946;
   wire v3_1517448501_947;
   wire v3_1517448501_948;
   wire v3_1517448501_949;
   wire v3_1517448501_950;
   wire v3_1517448501_951;
   wire v3_1517448501_952;
   wire v3_1517448501_953;
   wire v3_1517448501_954;
   wire v3_1517448501_955;
   wire f011;
   wire v3_1517448501_957;
   wire v3_1517448501_958;
   wire v3_1517448501_959;
   wire v3_1517448501_960;
   wire v3_1517448501_961;
   wire v3_1517448501_962;
   wire v3_1517448501_963;
   wire v3_1517448501_964;
   wire v3_1517448501_965;
   wire v3_1517448501_966;
   wire v3_1517448501_967;
   wire v3_1517448501_968;
   wire v3_1517448501_969;
   wire v3_1517448501_970;
   wire v3_1517448501_971;
   wire v3_1517448501_972;
   wire v3_1517448501_973;
   wire v3_1517448501_974;
   wire v3_1517448501_975;
   wire v3_1517448501_976;
   wire v3_1517448501_977;
   wire v3_1517448501_978;
   wire v3_1517448501_979;
   wire v3_1517448501_980;
   wire v3_1517448501_981;
   wire v3_1517448501_982;
   wire v3_1517448501_983;
   wire v3_1517448501_984;
   wire v3_1517448501_985;
   wire v3_1517448501_986;
   wire v3_1517448501_987;
   wire v3_1517448501_988;
   wire v3_1517448501_989;
   wire v3_1517448501_990;
   wire v3_1517448501_991;
   wire v3_1517448501_992;
   wire v3_1517448501_993;
   wire v3_1517448501_994;
   wire v3_1517448501_995;
   wire v3_1517448501_996;
   wire v3_1517448501_997;
   wire v3_1517448501_998;
   wire v3_1517448501_999;
   wire v3_1517448501_1000;
   wire v3_1517448501_1001;
   wire v3_1517448501_1002;
   wire v3_1517448501_1003;
   wire v3_1517448501_1004;
   wire v3_1517448501_1005;
   wire v3_1517448501_1006;
   wire v3_1517448501_1007;
   wire v3_1517448501_1008;
   wire v3_1517448501_1009;
   wire v3_1517448501_1010;
   wire v3_1517448501_1011;
   wire v3_1517448501_1012;
   wire v3_1517448501_1013;
   wire v3_1517448501_1014;
   wire v3_1517448501_1015;
   wire v3_1517448501_1016;
   wire v3_1517448501_1017;
   wire v3_1517448501_1018;
   wire v3_1517448501_1019;
   wire v3_1517448501_1020;
   wire v3_1517448501_1021;
   wire v3_1517448501_1022;
   wire v3_1517448501_1023;
   wire v3_1517448501_1024;
   wire v3_1517448501_1025;
   wire v3_1517448501_1026;
   wire f012;
   wire v3_1517448501_1028;
   wire f013;
   wire v3_1517448501_1030;
   wire v3_1517448501_1031;
   wire v3_1517448501_1032;
   wire v3_1517448501_1033;
   wire v3_1517448501_1034;
   wire v3_1517448501_1035;
   wire v3_1517448501_1036;
   wire v3_1517448501_1037;
   wire v3_1517448501_1038;
   wire v3_1517448501_1039;
   wire v3_1517448501_1040;
   wire v3_1517448501_1041;
   wire v3_1517448501_1042;
   wire v3_1517448501_1043;
   wire v3_1517448501_1044;
   wire v3_1517448501_1045;
   wire v3_1517448501_1046;
   wire v3_1517448501_1047;
   wire v3_1517448501_1048;
   wire v3_1517448501_1049;
   wire v3_1517448501_1050;
   wire v3_1517448501_1051;
   wire v3_1517448501_1052;
   wire v3_1517448501_1053;
   wire v3_1517448501_1054;
   wire v3_1517448501_1055;
   wire v3_1517448501_1056;
   wire v3_1517448501_1057;
   wire v3_1517448501_1058;
   wire v3_1517448501_1059;
   wire v3_1517448501_1060;
   wire v3_1517448501_1061;
   wire v3_1517448501_1062;
   wire v3_1517448501_1063;
   wire v3_1517448501_1064;
   wire v3_1517448501_1065;
   wire v3_1517448501_1066;
   wire v3_1517448501_1067;
   wire v3_1517448501_1068;
   wire v3_1517448501_1069;
   wire v3_1517448501_1070;
   wire v3_1517448501_1071;
   wire v3_1517448501_1072;
   wire v3_1517448501_1073;
   wire f015;
   wire v3_1517448501_1075;
   wire v3_1517448501_1076;
   wire v3_1517448501_1077;
   wire v3_1517448501_1078;
   wire v3_1517448501_1079;
   wire v3_1517448501_1080;
   wire v3_1517448501_1081;
   wire v3_1517448501_1082;
   wire v3_1517448501_1083;
   wire v3_1517448501_1084;
   wire v3_1517448501_1085;
   wire v3_1517448501_1086;
   wire v3_1517448501_1087;
   wire v3_1517448501_1088;
   wire v3_1517448501_1089;
   wire v3_1517448501_1090;
   wire v3_1517448501_1091;
   wire v3_1517448501_1092;
   wire v3_1517448501_1093;
   wire v3_1517448501_1094;
   wire v3_1517448501_1095;
   wire v3_1517448501_1096;
   wire v3_1517448501_1097;
   wire v3_1517448501_1098;
   wire v3_1517448501_1099;
   wire v3_1517448501_1100;
   wire v3_1517448501_1101;
   wire v3_1517448501_1102;
   wire v3_1517448501_1103;
   wire v3_1517448501_1104;
   wire v3_1517448501_1105;
   wire v3_1517448501_1106;
   wire v3_1517448501_1107;
   wire v3_1517448501_1108;
   wire v3_1517448501_1109;
   wire v3_1517448501_1110;
   wire v3_1517448501_1111;
   wire v3_1517448501_1112;
   wire v3_1517448501_1113;
   wire v3_1517448501_1114;
   wire v3_1517448501_1115;
   wire v3_1517448501_1116;
   wire v3_1517448501_1117;
   wire v3_1517448501_1118;
   wire v3_1517448501_1119;
   wire v3_1517448501_1120;
   wire v3_1517448501_1121;
   wire v3_1517448501_1122;
   wire v3_1517448501_1123;
   wire v3_1517448501_1124;
   wire v3_1517448501_1125;
   wire v3_1517448501_1126;
   wire v3_1517448501_1127;
   wire v3_1517448501_1128;
   wire v3_1517448501_1129;
   wire v3_1517448501_1130;
   wire v3_1517448501_1131;
   wire v3_1517448501_1132;
   wire v3_1517448501_1133;
   wire v3_1517448501_1134;
   wire v3_1517448501_1135;
   wire v3_1517448501_1136;
   wire v3_1517448501_1137;
   wire v3_1517448501_1138;
   wire v3_1517448501_1139;
   wire v3_1517448501_1140;
   wire v3_1517448501_1141;
   wire v3_1517448501_1142;
   wire v3_1517448501_1143;
   wire v3_1517448501_1144;
   wire f016;
   wire v3_1517448501_1146;
   wire f017;
   wire v3_1517448501_1148;
   wire v3_1517448501_1149;
   wire v3_1517448501_1150;
   wire v3_1517448501_1151;
   wire v3_1517448501_1152;
   wire v3_1517448501_1153;
   wire v3_1517448501_1154;
   wire v3_1517448501_1155;
   wire v3_1517448501_1156;
   wire v3_1517448501_1157;
   wire v3_1517448501_1158;
   wire v3_1517448501_1159;
   wire v3_1517448501_1160;
   wire v3_1517448501_1161;
   wire v3_1517448501_1162;
   wire v3_1517448501_1163;
   wire v3_1517448501_1164;
   wire v3_1517448501_1165;
   wire f018;
   wire v3_1517448501_1167;
   wire v3_1517448501_1168;
   wire v3_1517448501_1169;
   wire v3_1517448501_1170;
   wire f025;
   wire v3_1517448501_1172;
   wire v3_1517448501_1173;
   wire v3_1517448501_1174;
   wire v3_1517448501_1175;
   wire v3_1517448501_1176;
   wire v3_1517448501_1177;
   wire f028;
   wire v3_1517448501_1179;
   wire v3_1517448501_1180;
   wire v3_1517448501_1181;
   wire v3_1517448501_1182;
   wire v3_1517448501_1183;
   wire v3_1517448501_1184;
   wire f033;
   wire v3_1517448501_1186;
   wire v3_1517448501_1187;
   wire v3_1517448501_1188;
   wire v3_1517448501_1189;
   wire f035;
   wire v3_1517448501_1191;
   wire v3_1517448501_1192;
   wire v3_1517448501_1193;
   wire v3_1517448501_1194;
   wire v3_1517448501_1195;
   wire v3_1517448501_1196;
   wire v3_1517448501_1197;
   wire v3_1517448501_1198;
   wire v3_1517448501_1199;
   wire v3_1517448501_1200;
   wire v3_1517448501_1201;
   wire v3_1517448501_1202;
   wire v3_1517448501_1203;
   wire f019;
   wire v3_1517448501_1205;
   wire f020;
   wire v3_1517448501_1207;
   wire v3_1517448501_1208;
   wire v3_1517448501_1209;
   wire v3_1517448501_1210;
   wire v3_1517448501_1211;
   wire v3_1517448501_1212;
   wire v3_1517448501_1213;
   wire v3_1517448501_1214;
   wire v3_1517448501_1215;
   wire v3_1517448501_1216;
   wire v3_1517448501_1217;
   wire v3_1517448501_1218;
   wire v3_1517448501_1219;
   wire v3_1517448501_1220;
   wire v3_1517448501_1221;
   wire v3_1517448501_1222;
   wire v3_1517448501_1223;
   wire v3_1517448501_1224;
   wire f023;
   wire v3_1517448501_1226;
   wire v3_1517448501_1227;
   wire v3_1517448501_1228;
   wire v3_1517448501_1229;
   wire v3_1517448501_1230;
   wire v3_1517448501_1231;
   wire v3_1517448501_1232;
   wire v3_1517448501_1233;
   wire v3_1517448501_1234;
   wire v3_1517448501_1235;
   wire v3_1517448501_1236;
   wire v3_1517448501_1237;
   wire v3_1517448501_1238;
   wire v3_1517448501_1239;
   wire v3_1517448501_1240;
   wire v3_1517448501_1241;
   wire v3_1517448501_1242;
   wire f029;
   wire v3_1517448501_1244;
   wire f030;
   wire v3_1517448501_1246;
   wire v3_1517448501_1247;
   wire v3_1517448501_1248;
   wire v3_1517448501_1249;
   wire v3_1517448501_1250;
   wire v3_1517448501_1251;
   wire v3_1517448501_1252;
   wire v3_1517448501_1253;
   wire v3_1517448501_1254;
   wire v3_1517448501_1255;
   wire v3_1517448501_1256;
   wire v3_1517448501_1257;
   wire v3_1517448501_1258;
   wire v3_1517448501_1259;
   wire v3_1517448501_1260;
   wire v3_1517448501_1261;
   wire v3_1517448501_1262;
   wire v3_1517448501_1263;
   wire v3_1517448501_1264;
   wire [31:0] v3_1517448501_1265;
   wire [31:0] v3_1517448501_1266;
   wire v3_1517448501_1267;
   wire v3_1517448501_1268;
   wire [31:0] v3_1517448501_1269;
   wire [31:0] v3_1517448501_1270;
   wire [31:0] v3_1517448501_1271;
   wire [31:0] v3_1517448501_1272;
   wire [31:0] v3_1517448501_1273;
   wire [31:0] v3_1517448501_1274;
   wire [31:0] v3_1517448501_1275;
   wire v3_1517448501_1276;
   wire [31:0] v3_1517448501_1277;
   wire v3_1517448501_1278;
   wire v3_1517448501_1279;
   wire v3_1517448501_1280;
   wire [31:0] v3_1517448501_1281;
   wire [31:0] v3_1517448501_1282;
   wire [31:0] v3_1517448501_1283;
   wire [31:0] v3_1517448501_1284;
   wire [31:0] v3_1517448501_1285;
   wire [31:0] v3_1517448501_1286;
   wire [31:0] v3_1517448501_1287;
   wire v3_1517448501_1288;
   wire v3_1517448501_1289;
   wire v3_1517448501_1290;
   wire v3_1517448501_1291;
   wire v3_1517448501_1292;
   wire v3_1517448501_1293;
   wire v3_1517448501_1294;
   wire v3_1517448501_1295;
   wire v3_1517448501_1296;
   wire [31:0] v3_1517448501_1297;
   wire [31:0] v3_1517448501_1298;
   wire v3_1517448501_1299;
   wire v3_1517448501_1300;
   wire [31:0] v3_1517448501_1301;
   wire [31:0] v3_1517448501_1302;
   wire [31:0] v3_1517448501_1303;
   wire [31:0] v3_1517448501_1304;
   wire [31:0] v3_1517448501_1305;
   wire [31:0] v3_1517448501_1306;
   wire [31:0] v3_1517448501_1307;
   wire v3_1517448501_1308;
   wire [31:0] v3_1517448501_1309;
   wire [31:0] v3_1517448501_1310;
   wire v3_1517448501_1311;
   wire v3_1517448501_1312;
   wire v3_1517448501_1313;
   wire [31:0] v3_1517448501_1314;
   wire [31:0] v3_1517448501_1315;
   wire [31:0] v3_1517448501_1316;
   wire [31:0] v3_1517448501_1317;
   wire [31:0] v3_1517448501_1318;
   wire [31:0] v3_1517448501_1319;
   wire [31:0] v3_1517448501_1320;
   wire v3_1517448501_1321;
   wire v3_1517448501_1322;
   wire v3_1517448501_1323;
   wire v3_1517448501_1324;
   wire v3_1517448501_1325;
   wire v3_1517448501_1326;
   wire v3_1517448501_1327;
   wire v3_1517448501_1328;
   wire v3_1517448501_1329;
   wire v3_1517448501_1330;
   wire [31:0] v3_1517448501_1331;
   wire [31:0] v3_1517448501_1332;
   wire v3_1517448501_1333;
   wire v3_1517448501_1334;
   wire [31:0] v3_1517448501_1335;
   wire [31:0] v3_1517448501_1336;
   wire [31:0] v3_1517448501_1337;
   wire [31:0] v3_1517448501_1338;
   wire [31:0] v3_1517448501_1339;
   wire [31:0] v3_1517448501_1340;
   wire [31:0] v3_1517448501_1341;
   wire v3_1517448501_1342;
   wire [31:0] v3_1517448501_1343;
   wire [31:0] v3_1517448501_1344;
   wire v3_1517448501_1345;
   wire v3_1517448501_1346;
   wire v3_1517448501_1347;
   wire [31:0] v3_1517448501_1348;
   wire [31:0] v3_1517448501_1349;
   wire [31:0] v3_1517448501_1350;
   wire [31:0] v3_1517448501_1351;
   wire [31:0] v3_1517448501_1352;
   wire [31:0] v3_1517448501_1353;
   wire [31:0] v3_1517448501_1354;
   wire v3_1517448501_1355;
   wire v3_1517448501_1356;
   wire v3_1517448501_1357;
   wire v3_1517448501_1358;
   wire v3_1517448501_1359;
   wire v3_1517448501_1360;
   wire v3_1517448501_1361;
   wire v3_1517448501_1362;
   wire v3_1517448501_1363;
   wire v3_1517448501_1364;
   wire [31:0] v3_1517448501_1365;
   wire [31:0] v3_1517448501_1366;
   wire v3_1517448501_1367;
   wire v3_1517448501_1368;
   wire v3_1517448501_1369;
   wire [31:0] v3_1517448501_1370;
   wire [31:0] v3_1517448501_1371;
   wire [31:0] v3_1517448501_1372;
   wire [31:0] v3_1517448501_1373;
   wire [31:0] v3_1517448501_1374;
   wire [31:0] v3_1517448501_1375;
   wire [31:0] v3_1517448501_1376;
   wire v3_1517448501_1377;
   wire v3_1517448501_1378;
   wire v3_1517448501_1379;
   wire v3_1517448501_1380;
   wire v3_1517448501_1381;
   wire v3_1517448501_1382;
   wire v3_1517448501_1383;
   wire v3_1517448501_1384;
   wire v3_1517448501_1385;
   wire [31:0] v3_1517448501_1386;
   wire v3_1517448501_1387;
   wire v3_1517448501_1388;
   wire v3_1517448501_1389;
   wire v3_1517448501_1390;
   wire v3_1517448501_1391;
   wire v3_1517448501_1392;
   wire v3_1517448501_1393;
   wire v3_1517448501_1394;
   wire v3_1517448501_1395;
   wire v3_1517448501_1396;
   wire v3_1517448501_1397;
   wire [31:0] v3_1517448501_1398;
   wire [31:0] v3_1517448501_1399;
   wire v3_1517448501_1400;
   wire v3_1517448501_1401;
   wire v3_1517448501_1402;
   wire [31:0] v3_1517448501_1403;
   wire [31:0] v3_1517448501_1404;
   wire [31:0] v3_1517448501_1405;
   wire [31:0] v3_1517448501_1406;
   wire [31:0] v3_1517448501_1407;
   wire [31:0] v3_1517448501_1408;
   wire [31:0] v3_1517448501_1409;
   wire v3_1517448501_1410;
   wire v3_1517448501_1411;
   wire v3_1517448501_1412;
   wire v3_1517448501_1413;
   wire v3_1517448501_1414;
   wire v3_1517448501_1415;
   wire v3_1517448501_1416;
   wire v3_1517448501_1417;
   wire v3_1517448501_1418;
   wire [31:0] v3_1517448501_1419;
   wire v3_1517448501_1420;
   wire v3_1517448501_1421;
   wire v3_1517448501_1422;
   wire v3_1517448501_1423;
   wire v3_1517448501_1424;
   wire v3_1517448501_1425;
   wire v3_1517448501_1426;
   wire v3_1517448501_1427;
   wire v3_1517448501_1428;
   wire v3_1517448501_1429;
   wire v3_1517448501_1430;
   wire [31:0] v3_1517448501_1431;
   wire [31:0] v3_1517448501_1432;
   wire v3_1517448501_1433;
   wire v3_1517448501_1434;
   wire v3_1517448501_1435;
   wire [31:0] v3_1517448501_1436;
   wire [31:0] v3_1517448501_1437;
   wire [31:0] v3_1517448501_1438;
   wire [31:0] v3_1517448501_1439;
   wire [31:0] v3_1517448501_1440;
   wire [31:0] v3_1517448501_1441;
   wire [31:0] v3_1517448501_1442;
   wire v3_1517448501_1443;
   wire v3_1517448501_1444;
   wire v3_1517448501_1445;
   wire v3_1517448501_1446;
   wire v3_1517448501_1447;
   wire v3_1517448501_1448;
   wire v3_1517448501_1449;
   wire v3_1517448501_1450;
   wire v3_1517448501_1451;
   wire [31:0] v3_1517448501_1452;
   wire v3_1517448501_1453;
   wire v3_1517448501_1454;
   wire v3_1517448501_1455;
   wire v3_1517448501_1456;
   wire v3_1517448501_1457;
   wire v3_1517448501_1458;
   wire v3_1517448501_1459;
   wire v3_1517448501_1460;
   wire v3_1517448501_1461;
   wire v3_1517448501_1462;
   wire v3_1517448501_1463;
   wire v3_1517448501_1464;
   wire v3_1517448501_1465;
   wire v3_1517448501_1466;
   wire [31:0] v3_1517448501_1467;
   wire [31:0] v3_1517448501_1468;
   wire [31:0] v3_1517448501_1469;
   wire [31:0] v3_1517448501_1470;
   wire v3_1517448501_1471;
   wire [31:0] v3_1517448501_1472;
   wire v3_1517448501_1473;
   wire v3_1517448501_1474;
   wire v3_1517448501_1475;
   wire [31:0] v3_1517448501_1476;
   wire [31:0] v3_1517448501_1477;
   wire [31:0] v3_1517448501_1478;
   wire [31:0] v3_1517448501_1479;
   wire [31:0] v3_1517448501_1480;
   wire [31:0] v3_1517448501_1481;
   wire [31:0] v3_1517448501_1482;
   wire v3_1517448501_1483;
   wire v3_1517448501_1484;
   wire v3_1517448501_1485;
   wire v3_1517448501_1486;
   wire v3_1517448501_1487;
   wire v3_1517448501_1488;
   wire v3_1517448501_1489;
   wire v3_1517448501_1490;
   wire v3_1517448501_1491;
   wire [31:0] v3_1517448501_1492;
   wire v3_1517448501_1493;
   wire v3_1517448501_1494;
   wire [31:0] v3_1517448501_1495;
   wire [31:0] v3_1517448501_1496;
   wire [31:0] v3_1517448501_1497;
   wire [31:0] v3_1517448501_1498;
   wire [31:0] v3_1517448501_1499;
   wire [31:0] v3_1517448501_1500;
   wire [31:0] v3_1517448501_1501;
   wire v3_1517448501_1502;
   wire v3_1517448501_1503;
   wire v3_1517448501_1504;
   wire v3_1517448501_1505;
   wire v3_1517448501_1506;
   wire v3_1517448501_1507;
   wire v3_1517448501_1508;
   wire v3_1517448501_1509;
   wire v3_1517448501_1510;
   wire v3_1517448501_1511;
   wire v3_1517448501_1512;
   wire v3_1517448501_1513;
   wire v3_1517448501_1514;
   wire v3_1517448501_1515;
   wire v3_1517448501_1516;
   wire [31:0] v3_1517448501_1517;
   wire v3_1517448501_1518;
   wire v3_1517448501_1519;
   wire [31:0] v3_1517448501_1520;
   wire [31:0] v3_1517448501_1521;
   wire [31:0] v3_1517448501_1522;
   wire [31:0] v3_1517448501_1523;
   wire [31:0] v3_1517448501_1524;
   wire [31:0] v3_1517448501_1525;
   wire [31:0] v3_1517448501_1526;
   wire [31:0] v3_1517448501_1527;
   wire v3_1517448501_1528;
   wire v3_1517448501_1529;
   wire v3_1517448501_1530;
   wire [31:0] v3_1517448501_1531;
   wire [31:0] v3_1517448501_1532;
   wire [31:0] v3_1517448501_1533;
   wire [31:0] v3_1517448501_1534;
   wire [31:0] v3_1517448501_1535;
   wire [31:0] v3_1517448501_1536;
   wire [31:0] v3_1517448501_1537;
   wire v3_1517448501_1538;
   wire v3_1517448501_1539;
   wire v3_1517448501_1540;
   wire v3_1517448501_1541;
   wire v3_1517448501_1542;
   wire v3_1517448501_1543;
   wire v3_1517448501_1544;
   wire v3_1517448501_1545;
   wire v3_1517448501_1546;
   wire v3_1517448501_1547;
   wire v3_1517448501_1548;
   wire v3_1517448501_1549;
   wire v3_1517448501_1550;
   wire v3_1517448501_1551;
   wire v3_1517448501_1552;
   wire v3_1517448501_1553;
   wire v3_1517448501_1554;
   wire v3_1517448501_1555;
   wire v3_1517448501_1556;
   wire v3_1517448501_1557;
   wire v3_1517448501_1558;
   wire v3_1517448501_1559;
   wire v3_1517448501_1560;
   wire v3_1517448501_1561;
   wire v3_1517448501_1562;
   wire v3_1517448501_1563;
   wire v3_1517448501_1564;
   wire v3_1517448501_1565;
   wire v3_1517448501_1566;
   wire v3_1517448501_1567;
   wire v3_1517448501_1568;
   wire v3_1517448501_1569;
   wire v3_1517448501_1570;
   wire v3_1517448501_1571;
   wire v3_1517448501_1572;
   wire v3_1517448501_1573;
   wire v3_1517448501_1574;
   wire v3_1517448501_1575;
   wire v3_1517448501_1576;
   wire v3_1517448501_1577;
   wire v3_1517448501_1578;
   wire v3_1517448501_1579;
   wire v3_1517448501_1580;
   wire v3_1517448501_1581;
   wire v3_1517448501_1582;
   wire v3_1517448501_1583;
   wire v3_1517448501_1584;
   wire v3_1517448501_1585;
   wire v3_1517448501_1586;
   wire v3_1517448501_1587;
   wire v3_1517448501_1588;
   wire v3_1517448501_1589;
   wire v3_1517448501_1590;
   wire v3_1517448501_1591;
   wire v3_1517448501_1592;
   wire v3_1517448501_1593;
   wire v3_1517448501_1594;
   wire v3_1517448501_1595;
   wire v3_1517448501_1596;
   wire v3_1517448501_1597;
   wire v3_1517448501_1598;
   wire v3_1517448501_1599;
   wire v3_1517448501_1600;
   wire v3_1517448501_1601;
   wire v3_1517448501_1602;
   wire v3_1517448501_1603;
   wire v3_1517448501_1604;
   wire v3_1517448501_1605;
   wire v3_1517448501_1606;
   wire v3_1517448501_1607;
   wire v3_1517448501_1608;
   wire v3_1517448501_1609;
   wire v3_1517448501_1610;
   wire v3_1517448501_1611;
   wire v3_1517448501_1612;
   wire v3_1517448501_1613;
   wire v3_1517448501_1614;
   wire v3_1517448501_1615;
   wire v3_1517448501_1616;
   wire v3_1517448501_1617;
   wire v3_1517448501_1618;
   wire v3_1517448501_1619;
   wire v3_1517448501_1620;
   wire v3_1517448501_1621;
   wire v3_1517448501_1622;
   wire v3_1517448501_1623;
   wire v3_1517448501_1624;
   wire v3_1517448501_1625;
   wire v3_1517448501_1626;
   wire v3_1517448501_1627;
   wire v3_1517448501_1628;
   wire v3_1517448501_1629;
   wire v3_1517448501_1630;
   wire v3_1517448501_1631;
   wire v3_1517448501_1632;
   wire v3_1517448501_1633;
   wire v3_1517448501_1634;
   wire v3_1517448501_1635;
   wire v3_1517448501_1636;
   wire v3_1517448501_1637;
   wire v3_1517448501_1638;
   wire v3_1517448501_1639;
   wire v3_1517448501_1640;
   wire v3_1517448501_1641;
   wire v3_1517448501_1642;
   wire v3_1517448501_1643;
   wire v3_1517448501_1644;
   wire v3_1517448501_1645;
   wire v3_1517448501_1646;
   wire v3_1517448501_1647;
   wire v3_1517448501_1648;
   wire v3_1517448501_1649;
   wire v3_1517448501_1650;
   wire v3_1517448501_1651;
   wire v3_1517448501_1652;
   wire v3_1517448501_1653;
   wire v3_1517448501_1654;
   wire v3_1517448501_1655;
   wire v3_1517448501_1656;
   wire v3_1517448501_1657;
   wire v3_1517448501_1658;
   wire v3_1517448501_1659;
   wire v3_1517448501_1660;
   wire v3_1517448501_1661;
   wire v3_1517448501_1662;
   wire v3_1517448501_1663;
   wire v3_1517448501_1664;
   wire v3_1517448501_1665;
   wire v3_1517448501_1666;
   wire v3_1517448501_1667;
   wire v3_1517448501_1668;
   wire v3_1517448501_1669;
   wire v3_1517448501_1670;
   wire v3_1517448501_1671;
   wire v3_1517448501_1672;
   wire v3_1517448501_1673;
   wire v3_1517448501_1674;
   wire v3_1517448501_1675;
   wire v3_1517448501_1676;
   wire v3_1517448501_1677;
   wire v3_1517448501_1678;
   wire v3_1517448501_1679;
   wire v3_1517448501_1680;
   wire v3_1517448501_1681;
   wire v3_1517448501_1682;
   wire v3_1517448501_1683;
   wire v3_1517448501_1684;
   wire v3_1517448501_1685;
   wire v3_1517448501_1686;
   wire v3_1517448501_1687;
   wire v3_1517448501_1688;
   wire v3_1517448501_1689;
   wire v3_1517448501_1690;
   wire v3_1517448501_1691;
   wire v3_1517448501_1692;
   wire v3_1517448501_1693;
   wire v3_1517448501_1694;
   wire v3_1517448501_1695;
   wire v3_1517448501_1696;
   wire v3_1517448501_1697;
   wire v3_1517448501_1698;
   wire v3_1517448501_1699;
   wire v3_1517448501_1700;
   wire v3_1517448501_1701;
   wire v3_1517448501_1702;
   wire v3_1517448501_1703;
   wire v3_1517448501_1704;
   wire v3_1517448501_1705;
   wire v3_1517448501_1706;
   wire v3_1517448501_1707;
   wire v3_1517448501_1708;
   wire v3_1517448501_1709;
   wire v3_1517448501_1710;
   wire v3_1517448501_1711;
   wire v3_1517448501_1712;
   wire v3_1517448501_1713;
   wire v3_1517448501_1714;
   wire v3_1517448501_1715;
   wire v3_1517448501_1716;
   wire v3_1517448501_1717;
   wire v3_1517448501_1718;
   wire v3_1517448501_1719;
   wire v3_1517448501_1720;
   wire v3_1517448501_1721;
   wire v3_1517448501_1722;
   wire v3_1517448501_1723;
   wire v3_1517448501_1724;
   wire v3_1517448501_1725;
   wire v3_1517448501_1726;
   wire v3_1517448501_1727;
   wire v3_1517448501_1728;
   wire v3_1517448501_1729;
   wire v3_1517448501_1730;
   wire v3_1517448501_1731;
   wire v3_1517448501_1732;
   wire v3_1517448501_1733;
   wire v3_1517448501_1734;
   wire v3_1517448501_1735;
   wire v3_1517448501_1736;
   wire v3_1517448501_1737;
   wire v3_1517448501_1738;
   wire v3_1517448501_1739;
   wire v3_1517448501_1740;
   wire v3_1517448501_1741;
   wire v3_1517448501_1742;
   wire v3_1517448501_1743;
   wire v3_1517448501_1744;
   wire v3_1517448501_1745;
   wire v3_1517448501_1746;
   wire v3_1517448501_1747;
   wire v3_1517448501_1748;
   wire v3_1517448501_1749;
   wire v3_1517448501_1750;
   wire v3_1517448501_1751;
   wire v3_1517448501_1752;
   wire v3_1517448501_1753;
   wire v3_1517448501_1754;
   wire v3_1517448501_1755;
   wire v3_1517448501_1756;
   wire v3_1517448501_1757;
   wire v3_1517448501_1758;
   wire v3_1517448501_1759;
   wire v3_1517448501_1760;
   wire v3_1517448501_1761;
   wire v3_1517448501_1762;
   wire v3_1517448501_1763;
   wire v3_1517448501_1764;
   wire v3_1517448501_1765;
   wire v3_1517448501_1766;
   wire v3_1517448501_1767;
   wire v3_1517448501_1768;
   wire v3_1517448501_1769;
   wire v3_1517448501_1770;
   wire v3_1517448501_1771;
   wire v3_1517448501_1772;
   wire v3_1517448501_1773;
   wire v3_1517448501_1774;
   wire v3_1517448501_1775;
   wire v3_1517448501_1776;
   wire v3_1517448501_1777;
   wire v3_1517448501_1778;
   wire v3_1517448501_1779;
   wire v3_1517448501_1780;
   wire v3_1517448501_1781;
   wire v3_1517448501_1782;
   wire v3_1517448501_1783;
   wire v3_1517448501_1784;
   wire v3_1517448501_1785;
   wire v3_1517448501_1786;
   wire v3_1517448501_1787;
   wire v3_1517448501_1788;
   wire v3_1517448501_1789;
   wire [7:0] v3_1517448501_1790;
   wire v3_1517448501_1791;
   wire v3_1517448501_1792;
   wire v3_1517448501_1793;
   wire v3_1517448501_1794;
   wire v3_1517448501_1795;
   wire v3_1517448501_1796;
   wire v3_1517448501_1797;
   wire v3_1517448501_1798;
   wire v3_1517448501_1799;
   wire v3_1517448501_1800;
   wire v3_1517448501_1801;
   wire v3_1517448501_1802;
   wire v3_1517448501_1803;
   wire v3_1517448501_1804;
   wire v3_1517448501_1805;
   wire v3_1517448501_1806;
   wire v3_1517448501_1807;
   wire v3_1517448501_1808;
   wire v3_1517448501_1809;
   wire v3_1517448501_1810;
   wire v3_1517448501_1811;
   wire v3_1517448501_1812;
   wire v3_1517448501_1813;
   wire v3_1517448501_1814;
   wire v3_1517448501_1815;
   wire v3_1517448501_1816;
   wire v3_1517448501_1817;
   wire v3_1517448501_1818;
   wire v3_1517448501_1819;
   wire v3_1517448501_1820;
   wire v3_1517448501_1821;
   wire v3_1517448501_1822;
   wire v3_1517448501_1823;
   wire v3_1517448501_1824;
   wire v3_1517448501_1825;
   wire v3_1517448501_1826;
   wire v3_1517448501_1827;
   wire v3_1517448501_1828;
   wire v3_1517448501_1829;
   wire v3_1517448501_1830;
   wire v3_1517448501_1831;
   wire v3_1517448501_1832;
   wire v3_1517448501_1833;
   wire v3_1517448501_1834;
   wire v3_1517448501_1835;
   wire v3_1517448501_1836;
   wire v3_1517448501_1837;
   wire v3_1517448501_1838;
   wire v3_1517448501_1839;
   wire v3_1517448501_1840;
   wire v3_1517448501_1841;
   wire v3_1517448501_1842;
   wire v3_1517448501_1843;
   wire v3_1517448501_1844;
   wire v3_1517448501_1845;
   wire v3_1517448501_1846;
   wire v3_1517448501_1847;
   wire v3_1517448501_1848;
   wire v3_1517448501_1849;
   wire v3_1517448501_1850;
   wire v3_1517448501_1851;
   wire v3_1517448501_1852;
   wire v3_1517448501_1853;
   wire v3_1517448501_1854;
   wire v3_1517448501_1855;
   wire v3_1517448501_1856;
   wire v3_1517448501_1857;
   wire v3_1517448501_1858;
   wire v3_1517448501_1859;
   wire v3_1517448501_1860;
   wire v3_1517448501_1861;
   wire v3_1517448501_1862;
   wire v3_1517448501_1863;
   wire v3_1517448501_1864;
   wire v3_1517448501_1865;
   wire v3_1517448501_1866;
   wire v3_1517448501_1867;
   wire v3_1517448501_1868;
   wire v3_1517448501_1869;
   wire v3_1517448501_1870;
   wire v3_1517448501_1871;
   wire v3_1517448501_1872;
   wire v3_1517448501_1873;
   wire v3_1517448501_1874;
   wire v3_1517448501_1875;
   wire v3_1517448501_1876;
   wire v3_1517448501_1877;
   wire v3_1517448501_1878;
   wire v3_1517448501_1879;
   wire v3_1517448501_1880;
   wire v3_1517448501_1881;
   wire v3_1517448501_1882;
   wire v3_1517448501_1883;
   wire v3_1517448501_1884;
   wire v3_1517448501_1885;
   wire v3_1517448501_1886;
   wire v3_1517448501_1887;
   wire v3_1517448501_1888;
   wire v3_1517448501_1889;
   wire v3_1517448501_1890;
   wire v3_1517448501_1891;
   wire v3_1517448501_1892;
   wire v3_1517448501_1893;
   wire v3_1517448501_1894;
   wire v3_1517448501_1895;
   wire v3_1517448501_1896;
   wire v3_1517448501_1897;
   wire v3_1517448501_1898;
   wire v3_1517448501_1899;
   wire v3_1517448501_1900;
   wire v3_1517448501_1901;
   wire v3_1517448501_1902;
   wire v3_1517448501_1903;
   wire v3_1517448501_1904;
   wire v3_1517448501_1905;
   wire v3_1517448501_1906;
   wire v3_1517448501_1907;
   wire v3_1517448501_1908;
   wire v3_1517448501_1909;
   wire v3_1517448501_1910;
   wire v3_1517448501_1911;
   wire v3_1517448501_1912;
   wire v3_1517448501_1913;
   wire v3_1517448501_1914;
   wire v3_1517448501_1915;
   wire v3_1517448501_1916;
   wire v3_1517448501_1917;
   wire v3_1517448501_1918;
   wire v3_1517448501_1919;
   wire v3_1517448501_1920;
   wire v3_1517448501_1921;
   wire v3_1517448501_1922;
   wire v3_1517448501_1923;
   wire v3_1517448501_1924;
   wire v3_1517448501_1925;
   wire v3_1517448501_1926;
   wire v3_1517448501_1927;
   wire v3_1517448501_1928;
   wire v3_1517448501_1929;
   wire v3_1517448501_1930;
   wire v3_1517448501_1931;
   wire v3_1517448501_1932;
   wire v3_1517448501_1933;
   wire v3_1517448501_1934;
   wire v3_1517448501_1935;
   wire v3_1517448501_1936;
   wire v3_1517448501_1937;
   wire v3_1517448501_1938;
   wire v3_1517448501_1939;
   wire v3_1517448501_1940;
   wire v3_1517448501_1941;
   wire v3_1517448501_1942;
   wire v3_1517448501_1943;
   wire v3_1517448501_1944;
   wire v3_1517448501_1945;
   wire v3_1517448501_1946;
   wire v3_1517448501_1947;
   wire v3_1517448501_1948;
   wire v3_1517448501_1949;
   wire v3_1517448501_1950;
   wire v3_1517448501_1951;
   wire v3_1517448501_1952;
   wire v3_1517448501_1953;
   wire v3_1517448501_1954;
   wire v3_1517448501_1955;
   wire v3_1517448501_1956;
   wire v3_1517448501_1957;
   wire v3_1517448501_1958;
   wire v3_1517448501_1959;
   wire v3_1517448501_1960;
   wire v3_1517448501_1961;
   wire v3_1517448501_1962;
   wire v3_1517448501_1963;
   wire v3_1517448501_1964;
   wire v3_1517448501_1965;
   wire v3_1517448501_1966;
   wire v3_1517448501_1967;
   wire v3_1517448501_1968;
   wire v3_1517448501_1969;
   wire v3_1517448501_1970;
   wire v3_1517448501_1971;
   wire v3_1517448501_1972;
   wire v3_1517448501_1973;
   wire v3_1517448501_1974;
   wire v3_1517448501_1975;
   wire v3_1517448501_1976;
   wire v3_1517448501_1977;
   wire v3_1517448501_1978;
   wire v3_1517448501_1979;
   wire v3_1517448501_1980;
   wire v3_1517448501_1981;
   wire v3_1517448501_1982;
   wire v3_1517448501_1983;
   wire v3_1517448501_1984;
   wire v3_1517448501_1985;
   wire v3_1517448501_1986;
   wire v3_1517448501_1987;
   wire v3_1517448501_1988;
   wire v3_1517448501_1989;
   wire v3_1517448501_1990;
   wire v3_1517448501_1991;
   wire v3_1517448501_1992;
   wire v3_1517448501_1993;
   wire v3_1517448501_1994;
   wire v3_1517448501_1995;
   wire v3_1517448501_1996;
   wire v3_1517448501_1997;
   wire v3_1517448501_1998;
   wire v3_1517448501_1999;
   wire v3_1517448501_2000;
   wire v3_1517448501_2001;
   wire v3_1517448501_2002;
   wire v3_1517448501_2003;
   wire v3_1517448501_2004;
   wire v3_1517448501_2005;
   wire v3_1517448501_2006;
   wire v3_1517448501_2007;
   wire v3_1517448501_2008;
   wire v3_1517448501_2009;
   wire v3_1517448501_2010;
   wire v3_1517448501_2011;
   wire v3_1517448501_2012;
   wire v3_1517448501_2013;
   wire v3_1517448501_2014;
   wire v3_1517448501_2015;
   wire v3_1517448501_2016;
   wire v3_1517448501_2017;
   wire v3_1517448501_2018;
   wire v3_1517448501_2019;
   wire v3_1517448501_2020;
   wire v3_1517448501_2021;
   wire v3_1517448501_2022;
   wire v3_1517448501_2023;
   wire v3_1517448501_2024;
   wire v3_1517448501_2025;
   wire v3_1517448501_2026;
   wire v3_1517448501_2027;
   wire v3_1517448501_2028;
   wire v3_1517448501_2029;
   wire v3_1517448501_2030;
   wire v3_1517448501_2031;
   wire v3_1517448501_2032;
   wire v3_1517448501_2033;
   wire v3_1517448501_2034;
   wire v3_1517448501_2035;
   wire v3_1517448501_2036;
   wire v3_1517448501_2037;
   wire v3_1517448501_2038;
   wire v3_1517448501_2039;
   wire v3_1517448501_2040;
   wire v3_1517448501_2041;
   wire v3_1517448501_2042;
   wire v3_1517448501_2043;
   wire v3_1517448501_2044;
   wire v3_1517448501_2045;
   wire v3_1517448501_2046;
   wire v3_1517448501_2047;
   wire v3_1517448501_2048;
   wire v3_1517448501_2049;
   wire v3_1517448501_2050;
   wire v3_1517448501_2051;
   wire v3_1517448501_2052;
   wire v3_1517448501_2053;
   wire v3_1517448501_2054;
   wire v3_1517448501_2055;
   wire v3_1517448501_2056;
   wire v3_1517448501_2057;
   wire v3_1517448501_2058;
   wire v3_1517448501_2059;
   wire v3_1517448501_2060;
   wire v3_1517448501_2061;
   wire v3_1517448501_2062;
   wire v3_1517448501_2063;
   wire v3_1517448501_2064;
   wire v3_1517448501_2065;
   wire v3_1517448501_2066;
   wire v3_1517448501_2067;
   wire v3_1517448501_2068;
   wire v3_1517448501_2069;
   wire v3_1517448501_2070;
   wire v3_1517448501_2071;
   wire v3_1517448501_2072;
   wire v3_1517448501_2073;
   wire v3_1517448501_2074;
   wire v3_1517448501_2075;
   wire v3_1517448501_2076;
   wire v3_1517448501_2077;
   wire v3_1517448501_2078;
   wire v3_1517448501_2079;
   wire v3_1517448501_2080;
   wire v3_1517448501_2081;
   wire v3_1517448501_2082;
   wire v3_1517448501_2083;
   wire v3_1517448501_2084;
   wire v3_1517448501_2085;
   wire v3_1517448501_2086;
   wire v3_1517448501_2087;
   wire v3_1517448501_2088;
   wire v3_1517448501_2089;
   wire v3_1517448501_2090;
   wire v3_1517448501_2091;
   wire v3_1517448501_2092;
   wire v3_1517448501_2093;
   wire v3_1517448501_2094;
   wire v3_1517448501_2095;
   wire v3_1517448501_2096;
   wire v3_1517448501_2097;
   wire v3_1517448501_2098;
   wire v3_1517448501_2099;
   wire v3_1517448501_2100;
   wire v3_1517448501_2101;
   wire v3_1517448501_2102;
   wire v3_1517448501_2103;
   wire v3_1517448501_2104;
   wire v3_1517448501_2105;
   wire v3_1517448501_2106;
   wire v3_1517448501_2107;
   wire v3_1517448501_2108;
   wire v3_1517448501_2109;
   wire v3_1517448501_2110;
   wire v3_1517448501_2111;
   wire v3_1517448501_2112;
   wire v3_1517448501_2113;
   wire v3_1517448501_2114;
   wire v3_1517448501_2115;
   wire v3_1517448501_2116;
   wire v3_1517448501_2117;
   wire v3_1517448501_2118;
   wire v3_1517448501_2119;
   wire v3_1517448501_2120;
   wire v3_1517448501_2121;
   wire v3_1517448501_2122;
   wire v3_1517448501_2123;
   wire v3_1517448501_2124;
   wire v3_1517448501_2125;
   wire v3_1517448501_2126;
   wire v3_1517448501_2127;
   wire v3_1517448501_2128;
   wire v3_1517448501_2129;
   wire v3_1517448501_2130;
   wire v3_1517448501_2131;
   wire v3_1517448501_2132;
   wire v3_1517448501_2133;
   wire v3_1517448501_2134;
   wire v3_1517448501_2135;
   wire v3_1517448501_2136;
   wire v3_1517448501_2137;
   wire v3_1517448501_2138;
   wire v3_1517448501_2139;
   wire v3_1517448501_2140;
   wire v3_1517448501_2141;
   wire v3_1517448501_2142;
   wire v3_1517448501_2143;
   wire v3_1517448501_2144;
   wire v3_1517448501_2145;
   wire v3_1517448501_2146;
   wire v3_1517448501_2147;
   wire v3_1517448501_2148;
   wire v3_1517448501_2149;
   wire v3_1517448501_2150;
   wire v3_1517448501_2151;
   wire v3_1517448501_2152;
   wire v3_1517448501_2153;
   wire v3_1517448501_2154;
   wire v3_1517448501_2155;
   wire v3_1517448501_2156;
   wire v3_1517448501_2157;
   wire v3_1517448501_2158;
   wire v3_1517448501_2159;
   wire v3_1517448501_2160;
   wire v3_1517448501_2161;
   wire v3_1517448501_2162;
   wire v3_1517448501_2163;
   wire v3_1517448501_2164;
   wire v3_1517448501_2165;
   wire v3_1517448501_2166;
   wire v3_1517448501_2167;
   wire v3_1517448501_2168;
   wire v3_1517448501_2169;
   wire v3_1517448501_2170;
   wire v3_1517448501_2171;
   wire v3_1517448501_2172;
   wire v3_1517448501_2173;
   wire v3_1517448501_2174;
   wire v3_1517448501_2175;
   wire v3_1517448501_2176;
   wire v3_1517448501_2177;
   wire v3_1517448501_2178;
   wire v3_1517448501_2179;
   wire v3_1517448501_2180;
   wire v3_1517448501_2181;
   wire v3_1517448501_2182;
   wire v3_1517448501_2183;
   wire v3_1517448501_2184;
   wire v3_1517448501_2185;
   wire v3_1517448501_2186;
   wire v3_1517448501_2187;
   wire v3_1517448501_2188;
   wire v3_1517448501_2189;
   wire v3_1517448501_2190;
   wire v3_1517448501_2191;
   wire v3_1517448501_2192;
   wire v3_1517448501_2193;
   wire v3_1517448501_2194;
   wire v3_1517448501_2195;
   wire v3_1517448501_2196;
   wire v3_1517448501_2197;
   wire v3_1517448501_2198;
   wire v3_1517448501_2199;
   wire v3_1517448501_2200;
   wire v3_1517448501_2201;
   wire v3_1517448501_2202;
   wire v3_1517448501_2203;
   wire v3_1517448501_2204;
   wire v3_1517448501_2205;
   wire v3_1517448501_2206;
   wire v3_1517448501_2207;
   wire v3_1517448501_2208;
   wire v3_1517448501_2209;
   wire v3_1517448501_2210;
   wire v3_1517448501_2211;
   wire v3_1517448501_2212;
   wire v3_1517448501_2213;
   wire v3_1517448501_2214;
   wire v3_1517448501_2215;
   wire v3_1517448501_2216;
   wire v3_1517448501_2217;
   wire v3_1517448501_2218;
   wire v3_1517448501_2219;
   wire v3_1517448501_2220;
   wire v3_1517448501_2221;
   wire v3_1517448501_2222;
   wire v3_1517448501_2223;
   wire v3_1517448501_2224;
   wire v3_1517448501_2225;
   wire v3_1517448501_2226;
   wire v3_1517448501_2227;
   wire v3_1517448501_2228;
   wire v3_1517448501_2229;
   wire v3_1517448501_2230;
   wire v3_1517448501_2231;
   wire v3_1517448501_2232;
   wire v3_1517448501_2233;
   wire v3_1517448501_2234;
   wire v3_1517448501_2235;
   wire v3_1517448501_2236;
   wire v3_1517448501_2237;
   wire v3_1517448501_2238;
   wire v3_1517448501_2239;
   wire v3_1517448501_2240;
   wire v3_1517448501_2241;
   wire v3_1517448501_2242;
   wire v3_1517448501_2243;
   wire v3_1517448501_2244;
   wire v3_1517448501_2245;
   wire v3_1517448501_2246;
   wire v3_1517448501_2247;
   wire v3_1517448501_2248;
   wire v3_1517448501_2249;
   wire v3_1517448501_2250;
   wire v3_1517448501_2251;
   wire v3_1517448501_2252;
   wire v3_1517448501_2253;
   wire v3_1517448501_2254;
   wire v3_1517448501_2255;
   wire v3_1517448501_2256;
   wire v3_1517448501_2257;
   wire v3_1517448501_2258;
   wire v3_1517448501_2259;
   wire v3_1517448501_2260;
   wire v3_1517448501_2261;
   wire v3_1517448501_2262;
   wire v3_1517448501_2263;
   wire v3_1517448501_2264;
   wire v3_1517448501_2265;
   wire v3_1517448501_2266;
   wire v3_1517448501_2267;
   wire v3_1517448501_2268;
   wire v3_1517448501_2269;
   wire v3_1517448501_2270;
   wire v3_1517448501_2271;
   wire v3_1517448501_2272;
   wire v3_1517448501_2273;
   wire v3_1517448501_2274;
   wire v3_1517448501_2275;
   wire v3_1517448501_2276;
   wire v3_1517448501_2277;
   wire v3_1517448501_2278;
   wire v3_1517448501_2279;
   wire v3_1517448501_2280;
   wire v3_1517448501_2281;
   wire v3_1517448501_2282;
   wire v3_1517448501_2283;
   wire v3_1517448501_2284;
   wire v3_1517448501_2285;
   wire v3_1517448501_2286;
   wire v3_1517448501_2287;
   wire v3_1517448501_2288;
   wire v3_1517448501_2289;
   wire v3_1517448501_2290;
   wire v3_1517448501_2291;
   wire v3_1517448501_2292;
   wire v3_1517448501_2293;
   wire v3_1517448501_2294;
   wire v3_1517448501_2295;
   wire v3_1517448501_2296;
   wire v3_1517448501_2297;
   wire v3_1517448501_2298;
   wire v3_1517448501_2299;
   wire v3_1517448501_2300;
   wire v3_1517448501_2301;
   wire v3_1517448501_2302;
   wire v3_1517448501_2303;
   wire v3_1517448501_2304;
   wire v3_1517448501_2305;
   wire v3_1517448501_2306;
   wire v3_1517448501_2307;
   wire v3_1517448501_2308;
   wire v3_1517448501_2309;
   wire v3_1517448501_2310;
   wire v3_1517448501_2311;
   wire v3_1517448501_2312;
   wire v3_1517448501_2313;
   wire v3_1517448501_2314;
   wire v3_1517448501_2315;
   wire v3_1517448501_2316;
   wire v3_1517448501_2317;
   wire v3_1517448501_2318;
   wire v3_1517448501_2319;
   wire v3_1517448501_2320;
   wire v3_1517448501_2321;
   wire v3_1517448501_2322;
   wire v3_1517448501_2323;
   wire v3_1517448501_2324;
   wire v3_1517448501_2325;
   wire v3_1517448501_2326;
   wire v3_1517448501_2327;
   wire v3_1517448501_2328;
   wire v3_1517448501_2329;
   wire v3_1517448501_2330;
   wire v3_1517448501_2331;
   wire v3_1517448501_2332;
   wire v3_1517448501_2333;
   wire v3_1517448501_2334;
   wire v3_1517448501_2335;
   wire v3_1517448501_2336;
   wire v3_1517448501_2337;
   wire v3_1517448501_2338;
   wire v3_1517448501_2339;
   wire v3_1517448501_2340;
   wire v3_1517448501_2341;
   wire v3_1517448501_2342;
   wire v3_1517448501_2343;
   wire v3_1517448501_2344;
   wire v3_1517448501_2345;
   wire v3_1517448501_2346;
   wire v3_1517448501_2347;
   wire v3_1517448501_2348;
   wire v3_1517448501_2349;
   wire v3_1517448501_2350;
   wire v3_1517448501_2351;
   wire v3_1517448501_2352;
   wire v3_1517448501_2353;
   wire v3_1517448501_2354;
   wire v3_1517448501_2355;
   wire v3_1517448501_2356;
   wire v3_1517448501_2357;
   wire v3_1517448501_2358;
   wire v3_1517448501_2359;
   wire v3_1517448501_2360;
   wire v3_1517448501_2361;
   wire v3_1517448501_2362;
   wire v3_1517448501_2363;
   wire v3_1517448501_2364;
   wire v3_1517448501_2365;
   wire v3_1517448501_2366;
   wire v3_1517448501_2367;
   wire v3_1517448501_2368;
   wire v3_1517448501_2369;
   wire v3_1517448501_2370;
   wire v3_1517448501_2371;
   wire v3_1517448501_2372;
   wire v3_1517448501_2373;
   wire v3_1517448501_2374;
   wire v3_1517448501_2375;
   wire v3_1517448501_2376;
   wire v3_1517448501_2377;
   wire v3_1517448501_2378;
   wire v3_1517448501_2379;
   wire v3_1517448501_2380;
   wire v3_1517448501_2381;
   wire v3_1517448501_2382;
   wire v3_1517448501_2383;
   wire v3_1517448501_2384;
   wire v3_1517448501_2385;
   wire v3_1517448501_2386;
   wire v3_1517448501_2387;
   wire v3_1517448501_2388;
   wire v3_1517448501_2389;
   wire v3_1517448501_2390;
   wire v3_1517448501_2391;
   wire v3_1517448501_2392;
   wire v3_1517448501_2393;
   wire v3_1517448501_2394;
   wire v3_1517448501_2395;
   wire v3_1517448501_2396;
   wire v3_1517448501_2397;
   wire v3_1517448501_2398;
   wire v3_1517448501_2399;
   wire v3_1517448501_2400;
   wire v3_1517448501_2401;
   wire v3_1517448501_2402;
   wire v3_1517448501_2403;
   wire v3_1517448501_2404;
   wire v3_1517448501_2405;
   wire v3_1517448501_2406;
   wire v3_1517448501_2407;
   wire v3_1517448501_2408;
   wire v3_1517448501_2409;
   wire v3_1517448501_2410;
   wire v3_1517448501_2411;
   wire v3_1517448501_2412;
   wire v3_1517448501_2413;
   wire v3_1517448501_2414;
   wire v3_1517448501_2415;
   wire v3_1517448501_2416;
   wire v3_1517448501_2417;
   wire v3_1517448501_2418;
   wire v3_1517448501_2419;
   wire v3_1517448501_2420;
   wire v3_1517448501_2421;
   wire v3_1517448501_2422;
   wire v3_1517448501_2423;
   wire v3_1517448501_2424;
   wire v3_1517448501_2425;
   wire v3_1517448501_2426;
   wire v3_1517448501_2427;
   wire v3_1517448501_2428;
   wire v3_1517448501_2429;
   wire v3_1517448501_2430;
   wire v3_1517448501_2431;
   wire v3_1517448501_2432;
   wire v3_1517448501_2433;
   wire v3_1517448501_2434;
   wire v3_1517448501_2435;
   wire v3_1517448501_2436;
   wire v3_1517448501_2437;
   wire v3_1517448501_2438;
   wire v3_1517448501_2439;
   wire v3_1517448501_2440;
   wire v3_1517448501_2441;
   wire v3_1517448501_2442;
   wire v3_1517448501_2443;
   wire v3_1517448501_2444;
   wire v3_1517448501_2445;
   wire v3_1517448501_2446;
   wire v3_1517448501_2447;
   wire v3_1517448501_2448;
   wire v3_1517448501_2449;
   wire v3_1517448501_2450;
   wire v3_1517448501_2451;
   wire v3_1517448501_2452;
   wire v3_1517448501_2453;
   wire v3_1517448501_2454;
   wire v3_1517448501_2455;
   wire v3_1517448501_2456;
   wire v3_1517448501_2457;
   wire v3_1517448501_2458;
   wire v3_1517448501_2459;
   wire v3_1517448501_2460;
   wire v3_1517448501_2461;
   wire v3_1517448501_2462;
   wire v3_1517448501_2463;
   wire v3_1517448501_2464;
   wire v3_1517448501_2465;
   wire v3_1517448501_2466;
   wire v3_1517448501_2467;
   wire v3_1517448501_2468;
   wire v3_1517448501_2469;
   wire v3_1517448501_2470;
   wire v3_1517448501_2471;
   wire v3_1517448501_2472;
   wire v3_1517448501_2473;
   wire v3_1517448501_2474;
   wire v3_1517448501_2475;
   wire v3_1517448501_2476;
   wire v3_1517448501_2477;
   wire v3_1517448501_2478;
   wire v3_1517448501_2479;
   wire v3_1517448501_2480;
   wire v3_1517448501_2481;
   wire v3_1517448501_2482;
   wire v3_1517448501_2483;
   wire v3_1517448501_2484;
   wire v3_1517448501_2485;
   wire v3_1517448501_2486;
   wire v3_1517448501_2487;
   wire v3_1517448501_2488;
   wire v3_1517448501_2489;
   wire v3_1517448501_2490;
   wire v3_1517448501_2491;
   wire v3_1517448501_2492;
   wire v3_1517448501_2493;
   wire v3_1517448501_2494;
   wire v3_1517448501_2495;
   wire v3_1517448501_2496;
   wire v3_1517448501_2497;
   wire v3_1517448501_2498;
   wire v3_1517448501_2499;
   wire v3_1517448501_2500;
   wire v3_1517448501_2501;
   wire v3_1517448501_2502;
   wire v3_1517448501_2503;
   wire v3_1517448501_2504;
   wire v3_1517448501_2505;
   wire v3_1517448501_2506;
   wire v3_1517448501_2507;
   wire v3_1517448501_2508;
   wire v3_1517448501_2509;
   wire v3_1517448501_2510;
   wire v3_1517448501_2511;
   wire v3_1517448501_2512;
   wire v3_1517448501_2513;
   wire v3_1517448501_2514;
   wire v3_1517448501_2515;
   wire v3_1517448501_2516;
   wire v3_1517448501_2517;
   wire v3_1517448501_2518;
   wire v3_1517448501_2519;
   wire v3_1517448501_2520;
   wire v3_1517448501_2521;
   wire v3_1517448501_2522;
   wire v3_1517448501_2523;
   wire v3_1517448501_2524;
   wire v3_1517448501_2525;
   wire v3_1517448501_2526;
   wire v3_1517448501_2527;
   wire v3_1517448501_2528;
   wire v3_1517448501_2529;
   wire v3_1517448501_2530;
   wire v3_1517448501_2531;
   wire v3_1517448501_2532;
   wire v3_1517448501_2533;
   wire v3_1517448501_2534;
   wire v3_1517448501_2535;
   wire v3_1517448501_2536;
   wire v3_1517448501_2537;
   wire v3_1517448501_2538;
   wire v3_1517448501_2539;
   wire v3_1517448501_2540;
   wire v3_1517448501_2541;
   wire v3_1517448501_2542;
   wire v3_1517448501_2543;
   wire v3_1517448501_2544;
   wire v3_1517448501_2545;
   wire v3_1517448501_2546;
   wire v3_1517448501_2547;
   wire v3_1517448501_2548;
   wire v3_1517448501_2549;
   wire v3_1517448501_2550;
   wire v3_1517448501_2551;
   wire v3_1517448501_2552;
   wire v3_1517448501_2553;
   wire v3_1517448501_2554;
   wire v3_1517448501_2555;
   wire v3_1517448501_2556;
   wire v3_1517448501_2557;
   wire v3_1517448501_2558;
   wire v3_1517448501_2559;
   wire v3_1517448501_2560;
   wire v3_1517448501_2561;
   wire v3_1517448501_2562;
   wire v3_1517448501_2563;
   wire v3_1517448501_2564;
   wire v3_1517448501_2565;
   wire v3_1517448501_2566;
   wire v3_1517448501_2567;
   wire v3_1517448501_2568;
   wire v3_1517448501_2569;
   wire v3_1517448501_2570;
   wire v3_1517448501_2571;
   wire v3_1517448501_2572;
   wire v3_1517448501_2573;
   wire v3_1517448501_2574;
   wire v3_1517448501_2575;
   wire v3_1517448501_2576;
   wire v3_1517448501_2577;
   wire v3_1517448501_2578;
   wire v3_1517448501_2579;
   wire v3_1517448501_2580;
   wire v3_1517448501_2581;
   wire v3_1517448501_2582;
   wire v3_1517448501_2583;
   wire v3_1517448501_2584;
   wire v3_1517448501_2585;
   wire v3_1517448501_2586;
   wire v3_1517448501_2587;
   wire v3_1517448501_2588;
   wire v3_1517448501_2589;
   wire v3_1517448501_2590;
   wire v3_1517448501_2591;
   wire v3_1517448501_2592;
   wire v3_1517448501_2593;
   wire v3_1517448501_2594;
   wire v3_1517448501_2595;
   wire v3_1517448501_2596;
   wire v3_1517448501_2597;
   wire v3_1517448501_2598;
   wire v3_1517448501_2599;
   wire v3_1517448501_2600;
   wire v3_1517448501_2601;
   wire v3_1517448501_2602;
   wire v3_1517448501_2603;
   wire v3_1517448501_2604;
   wire v3_1517448501_2605;
   wire v3_1517448501_2606;
   wire v3_1517448501_2607;
   wire v3_1517448501_2608;
   wire v3_1517448501_2609;
   wire v3_1517448501_2610;
   wire v3_1517448501_2611;
   wire v3_1517448501_2612;
   wire v3_1517448501_2613;
   wire v3_1517448501_2614;
   wire v3_1517448501_2615;
   wire v3_1517448501_2616;
   wire v3_1517448501_2617;
   wire v3_1517448501_2618;
   wire v3_1517448501_2619;
   wire v3_1517448501_2620;
   wire v3_1517448501_2621;
   wire v3_1517448501_2622;
   wire v3_1517448501_2623;
   wire v3_1517448501_2624;
   wire v3_1517448501_2625;
   wire v3_1517448501_2626;
   wire v3_1517448501_2627;
   wire v3_1517448501_2628;
   wire v3_1517448501_2629;
   wire v3_1517448501_2630;
   wire v3_1517448501_2631;
   wire v3_1517448501_2632;
   wire v3_1517448501_2633;
   wire v3_1517448501_2634;
   wire v3_1517448501_2635;
   wire v3_1517448501_2636;
   wire v3_1517448501_2637;
   wire v3_1517448501_2638;
   wire v3_1517448501_2639;
   wire v3_1517448501_2640;
   wire v3_1517448501_2641;
   wire v3_1517448501_2642;
   wire v3_1517448501_2643;
   wire v3_1517448501_2644;
   wire v3_1517448501_2645;
   wire v3_1517448501_2646;
   wire v3_1517448501_2647;
   wire v3_1517448501_2648;
   wire v3_1517448501_2649;
   wire v3_1517448501_2650;
   wire v3_1517448501_2651;
   wire v3_1517448501_2652;
   wire v3_1517448501_2653;
   wire v3_1517448501_2654;
   wire v3_1517448501_2655;
   wire v3_1517448501_2656;
   wire v3_1517448501_2657;
   wire v3_1517448501_2658;
   wire v3_1517448501_2659;
   wire v3_1517448501_2660;
   wire v3_1517448501_2661;
   wire v3_1517448501_2662;
   wire v3_1517448501_2663;
   wire v3_1517448501_2664;
   wire v3_1517448501_2665;
   wire v3_1517448501_2666;
   wire v3_1517448501_2667;
   wire v3_1517448501_2668;
   wire v3_1517448501_2669;
   wire v3_1517448501_2670;
   wire v3_1517448501_2671;
   wire v3_1517448501_2672;
   wire v3_1517448501_2673;
   wire v3_1517448501_2674;
   wire v3_1517448501_2675;
   wire v3_1517448501_2676;
   wire v3_1517448501_2677;
   wire v3_1517448501_2678;
   wire v3_1517448501_2679;
   wire v3_1517448501_2680;
   wire v3_1517448501_2681;
   wire v3_1517448501_2682;
   wire v3_1517448501_2683;
   wire v3_1517448501_2684;
   wire v3_1517448501_2685;
   wire v3_1517448501_2686;
   wire v3_1517448501_2687;
   wire v3_1517448501_2688;
   wire v3_1517448501_2689;
   wire v3_1517448501_2690;
   wire v3_1517448501_2691;
   wire v3_1517448501_2692;
   wire v3_1517448501_2693;
   wire v3_1517448501_2694;
   wire v3_1517448501_2695;
   wire v3_1517448501_2696;
   wire v3_1517448501_2697;
   wire v3_1517448501_2698;
   wire v3_1517448501_2699;
   wire v3_1517448501_2700;
   wire v3_1517448501_2701;
   wire v3_1517448501_2702;
   wire v3_1517448501_2703;
   wire v3_1517448501_2704;
   wire v3_1517448501_2705;
   wire v3_1517448501_2706;
   wire v3_1517448501_2707;
   wire v3_1517448501_2708;
   wire v3_1517448501_2709;
   wire v3_1517448501_2710;
   wire v3_1517448501_2711;
   wire v3_1517448501_2712;
   wire v3_1517448501_2713;
   wire v3_1517448501_2714;
   wire v3_1517448501_2715;
   wire v3_1517448501_2716;
   wire v3_1517448501_2717;
   wire v3_1517448501_2718;
   wire v3_1517448501_2719;
   wire v3_1517448501_2720;
   wire v3_1517448501_2721;
   wire v3_1517448501_2722;
   wire v3_1517448501_2723;
   wire v3_1517448501_2724;
   wire v3_1517448501_2725;
   wire v3_1517448501_2726;
   wire v3_1517448501_2727;
   wire v3_1517448501_2728;
   wire v3_1517448501_2729;
   wire v3_1517448501_2730;
   wire v3_1517448501_2731;
   wire v3_1517448501_2732;
   wire v3_1517448501_2733;
   wire v3_1517448501_2734;
   wire v3_1517448501_2735;
   wire v3_1517448501_2736;
   wire v3_1517448501_2737;
   wire v3_1517448501_2738;
   wire v3_1517448501_2739;
   wire v3_1517448501_2740;
   wire v3_1517448501_2741;
   wire v3_1517448501_2742;
   wire v3_1517448501_2743;
   wire v3_1517448501_2744;
   wire v3_1517448501_2745;
   wire v3_1517448501_2746;
   wire v3_1517448501_2747;
   wire v3_1517448501_2748;
   wire v3_1517448501_2749;
   wire v3_1517448501_2750;
   wire v3_1517448501_2751;
   wire v3_1517448501_2752;
   wire v3_1517448501_2753;
   wire v3_1517448501_2754;
   wire v3_1517448501_2755;
   wire v3_1517448501_2756;
   wire v3_1517448501_2757;
   wire v3_1517448501_2758;
   wire v3_1517448501_2759;
   wire v3_1517448501_2760;
   wire v3_1517448501_2761;
   wire v3_1517448501_2762;
   wire v3_1517448501_2763;
   wire v3_1517448501_2764;
   wire v3_1517448501_2765;
   wire v3_1517448501_2766;
   wire v3_1517448501_2767;
   wire v3_1517448501_2768;
   wire v3_1517448501_2769;
   wire v3_1517448501_2770;
   wire v3_1517448501_2771;
   wire v3_1517448501_2772;
   wire v3_1517448501_2773;
   wire v3_1517448501_2774;
   wire v3_1517448501_2775;
   wire v3_1517448501_2776;
   wire v3_1517448501_2777;
   wire v3_1517448501_2778;
   wire v3_1517448501_2779;
   wire v3_1517448501_2780;
   wire v3_1517448501_2781;
   wire v3_1517448501_2782;
   wire v3_1517448501_2783;
   wire v3_1517448501_2784;
   wire v3_1517448501_2785;
   wire v3_1517448501_2786;
   wire v3_1517448501_2787;
   wire v3_1517448501_2788;
   wire v3_1517448501_2789;
   wire v3_1517448501_2790;
   wire v3_1517448501_2791;
   wire v3_1517448501_2792;
   wire v3_1517448501_2793;
   wire v3_1517448501_2794;
   wire v3_1517448501_2795;
   wire v3_1517448501_2796;
   wire v3_1517448501_2797;
   wire v3_1517448501_2798;
   wire v3_1517448501_2799;
   wire v3_1517448501_2800;
   wire v3_1517448501_2801;
   wire v3_1517448501_2802;
   wire v3_1517448501_2803;
   wire v3_1517448501_2804;
   wire v3_1517448501_2805;
   wire v3_1517448501_2806;
   wire v3_1517448501_2807;
   wire v3_1517448501_2808;
   wire v3_1517448501_2809;
   wire v3_1517448501_2810;
   wire v3_1517448501_2811;
   wire v3_1517448501_2812;
   wire v3_1517448501_2813;
   wire v3_1517448501_2814;
   wire v3_1517448501_2815;
   wire v3_1517448501_2816;
   wire v3_1517448501_2817;
   wire v3_1517448501_2818;
   wire v3_1517448501_2819;
   wire v3_1517448501_2820;
   wire v3_1517448501_2821;
   wire v3_1517448501_2822;
   wire v3_1517448501_2823;
   wire v3_1517448501_2824;
   wire v3_1517448501_2825;
   wire v3_1517448501_2826;
   wire v3_1517448501_2827;
   wire v3_1517448501_2828;
   wire v3_1517448501_2829;
   wire v3_1517448501_2830;
   wire v3_1517448501_2831;
   wire v3_1517448501_2832;
   wire v3_1517448501_2833;
   wire v3_1517448501_2834;
   wire v3_1517448501_2835;
   wire v3_1517448501_2836;
   wire v3_1517448501_2837;
   wire v3_1517448501_2838;
   wire v3_1517448501_2839;
   wire v3_1517448501_2840;
   wire v3_1517448501_2841;
   wire v3_1517448501_2842;
   wire v3_1517448501_2843;
   wire v3_1517448501_2844;
   wire v3_1517448501_2845;
   wire v3_1517448501_2846;
   wire v3_1517448501_2847;
   wire v3_1517448501_2848;
   wire v3_1517448501_2849;
   wire v3_1517448501_2850;
   wire v3_1517448501_2851;
   wire v3_1517448501_2852;
   wire v3_1517448501_2853;
   wire v3_1517448501_2854;
   wire v3_1517448501_2855;
   wire v3_1517448501_2856;
   wire v3_1517448501_2857;
   wire v3_1517448501_2858;
   wire v3_1517448501_2859;
   wire v3_1517448501_2860;
   wire v3_1517448501_2861;
   wire v3_1517448501_2862;
   wire v3_1517448501_2863;
   wire v3_1517448501_2864;
   wire v3_1517448501_2865;
   wire v3_1517448501_2866;
   wire v3_1517448501_2867;
   wire v3_1517448501_2868;
   wire v3_1517448501_2869;
   wire v3_1517448501_2870;
   wire v3_1517448501_2871;
   wire v3_1517448501_2872;
   wire v3_1517448501_2873;
   wire v3_1517448501_2874;
   wire v3_1517448501_2875;
   wire v3_1517448501_2876;
   wire v3_1517448501_2877;
   wire v3_1517448501_2878;
   wire v3_1517448501_2879;
   wire v3_1517448501_2880;
   wire v3_1517448501_2881;
   wire v3_1517448501_2882;
   wire v3_1517448501_2883;
   wire v3_1517448501_2884;
   wire v3_1517448501_2885;
   wire v3_1517448501_2886;
   wire v3_1517448501_2887;
   wire v3_1517448501_2888;
   wire v3_1517448501_2889;
   wire v3_1517448501_2890;
   wire v3_1517448501_2891;
   wire v3_1517448501_2892;
   wire v3_1517448501_2893;
   wire v3_1517448501_2894;
   wire v3_1517448501_2895;
   wire v3_1517448501_2896;
   wire v3_1517448501_2897;
   wire v3_1517448501_2898;
   wire v3_1517448501_2899;
   wire v3_1517448501_2900;
   wire v3_1517448501_2901;
   wire v3_1517448501_2902;
   wire v3_1517448501_2903;
   wire v3_1517448501_2904;
   wire v3_1517448501_2905;
   wire v3_1517448501_2906;
   wire v3_1517448501_2907;
   wire v3_1517448501_2908;
   wire v3_1517448501_2909;
   wire v3_1517448501_2910;
   wire v3_1517448501_2911;
   wire v3_1517448501_2912;
   wire v3_1517448501_2913;
   wire v3_1517448501_2914;
   wire v3_1517448501_2915;
   wire v3_1517448501_2916;
   wire v3_1517448501_2917;
   wire v3_1517448501_2918;
   wire v3_1517448501_2919;
   wire v3_1517448501_2920;
   wire v3_1517448501_2921;
   wire v3_1517448501_2922;
   wire v3_1517448501_2923;
   wire v3_1517448501_2924;
   wire v3_1517448501_2925;
   wire v3_1517448501_2926;
   wire v3_1517448501_2927;
   wire v3_1517448501_2928;
   wire v3_1517448501_2929;
   wire v3_1517448501_2930;
   wire v3_1517448501_2931;
   wire v3_1517448501_2932;
   wire v3_1517448501_2933;
   wire v3_1517448501_2934;
   wire v3_1517448501_2935;
   wire v3_1517448501_2936;
   wire v3_1517448501_2937;
   wire v3_1517448501_2938;
   wire v3_1517448501_2939;
   wire v3_1517448501_2940;
   wire v3_1517448501_2941;
   wire v3_1517448501_2942;
   wire v3_1517448501_2943;
   wire v3_1517448501_2944;
   wire v3_1517448501_2945;
   wire v3_1517448501_2946;
   wire v3_1517448501_2947;
   wire v3_1517448501_2948;
   wire v3_1517448501_2949;
   wire v3_1517448501_2950;
   wire v3_1517448501_2951;
   wire v3_1517448501_2952;
   wire v3_1517448501_2953;
   wire v3_1517448501_2954;
   wire v3_1517448501_2955;
   wire v3_1517448501_2956;
   wire v3_1517448501_2957;
   wire v3_1517448501_2958;
   wire v3_1517448501_2959;
   wire v3_1517448501_2960;
   wire v3_1517448501_2961;
   wire v3_1517448501_2962;
   wire v3_1517448501_2963;
   wire v3_1517448501_2964;
   wire v3_1517448501_2965;
   wire v3_1517448501_2966;
   wire v3_1517448501_2967;
   wire v3_1517448501_2968;
   wire v3_1517448501_2969;
   wire v3_1517448501_2970;
   wire v3_1517448501_2971;
   wire v3_1517448501_2972;
   wire v3_1517448501_2973;
   wire v3_1517448501_2974;
   wire v3_1517448501_2975;
   wire v3_1517448501_2976;
   wire v3_1517448501_2977;
   wire v3_1517448501_2978;
   wire v3_1517448501_2979;
   wire v3_1517448501_2980;
   wire v3_1517448501_2981;
   wire v3_1517448501_2982;
   wire v3_1517448501_2983;
   wire v3_1517448501_2984;
   wire v3_1517448501_2985;
   wire v3_1517448501_2986;
   wire v3_1517448501_2987;
   wire v3_1517448501_2988;
   wire v3_1517448501_2989;
   wire v3_1517448501_2990;
   wire v3_1517448501_2991;
   wire v3_1517448501_2992;
   wire v3_1517448501_2993;
   wire v3_1517448501_2994;
   wire v3_1517448501_2995;
   wire v3_1517448501_2996;
   wire v3_1517448501_2997;
   wire v3_1517448501_2998;
   wire v3_1517448501_2999;
   wire v3_1517448501_3000;
   wire v3_1517448501_3001;
   wire v3_1517448501_3002;
   wire v3_1517448501_3003;
   wire v3_1517448501_3004;
   wire v3_1517448501_3005;
   wire v3_1517448501_3006;
   wire v3_1517448501_3007;
   wire v3_1517448501_3008;
   wire v3_1517448501_3009;
   wire v3_1517448501_3010;
   wire v3_1517448501_3011;
   wire v3_1517448501_3012;
   wire v3_1517448501_3013;
   wire v3_1517448501_3014;
   wire v3_1517448501_3015;
   wire v3_1517448501_3016;
   wire v3_1517448501_3017;
   wire v3_1517448501_3018;
   wire v3_1517448501_3019;
   wire v3_1517448501_3020;
   wire v3_1517448501_3021;
   wire v3_1517448501_3022;
   wire v3_1517448501_3023;
   wire v3_1517448501_3024;
   wire v3_1517448501_3025;
   wire v3_1517448501_3026;
   wire v3_1517448501_3027;
   wire v3_1517448501_3028;
   wire v3_1517448501_3029;
   wire v3_1517448501_3030;
   wire v3_1517448501_3031;
   wire v3_1517448501_3032;
   wire v3_1517448501_3033;
   wire v3_1517448501_3034;
   wire v3_1517448501_3035;
   wire v3_1517448501_3036;
   wire v3_1517448501_3037;
   wire v3_1517448501_3038;
   wire v3_1517448501_3039;
   wire v3_1517448501_3040;
   wire v3_1517448501_3041;
   wire v3_1517448501_3042;
   wire v3_1517448501_3043;
   wire v3_1517448501_3044;
   wire v3_1517448501_3045;
   wire v3_1517448501_3046;
   wire v3_1517448501_3047;
   wire v3_1517448501_3048;
   wire v3_1517448501_3049;
   wire v3_1517448501_3050;
   wire v3_1517448501_3051;
   wire v3_1517448501_3052;
   wire v3_1517448501_3053;
   wire v3_1517448501_3054;
   wire v3_1517448501_3055;
   wire v3_1517448501_3056;
   wire v3_1517448501_3057;
   wire v3_1517448501_3058;
   wire v3_1517448501_3059;
   wire v3_1517448501_3060;
   wire v3_1517448501_3061;
   wire v3_1517448501_3062;
   wire v3_1517448501_3063;
   wire v3_1517448501_3064;
   wire v3_1517448501_3065;
   wire v3_1517448501_3066;
   wire v3_1517448501_3067;
   wire v3_1517448501_3068;
   wire v3_1517448501_3069;
   wire v3_1517448501_3070;
   wire v3_1517448501_3071;
   wire v3_1517448501_3072;
   wire v3_1517448501_3073;
   wire v3_1517448501_3074;
   wire v3_1517448501_3075;
   wire v3_1517448501_3076;
   wire v3_1517448501_3077;
   wire v3_1517448501_3078;
   wire v3_1517448501_3079;
   wire v3_1517448501_3080;
   wire v3_1517448501_3081;
   wire v3_1517448501_3082;
   wire v3_1517448501_3083;
   wire v3_1517448501_3084;
   wire v3_1517448501_3085;
   wire v3_1517448501_3086;
   wire v3_1517448501_3087;
   wire v3_1517448501_3088;
   wire v3_1517448501_3089;
   wire v3_1517448501_3090;
   wire v3_1517448501_3091;
   wire v3_1517448501_3092;
   wire v3_1517448501_3093;
   wire v3_1517448501_3094;
   wire v3_1517448501_3095;
   wire v3_1517448501_3096;
   wire v3_1517448501_3097;
   wire v3_1517448501_3098;
   wire v3_1517448501_3099;
   wire v3_1517448501_3100;
   wire v3_1517448501_3101;
   wire v3_1517448501_3102;
   wire v3_1517448501_3103;
   wire v3_1517448501_3104;
   wire v3_1517448501_3105;
   wire v3_1517448501_3106;
   wire v3_1517448501_3107;
   wire v3_1517448501_3108;
   wire v3_1517448501_3109;
   wire v3_1517448501_3110;
   wire v3_1517448501_3111;
   wire v3_1517448501_3112;
   wire v3_1517448501_3113;
   wire v3_1517448501_3114;
   wire v3_1517448501_3115;
   wire v3_1517448501_3116;
   wire v3_1517448501_3117;
   wire v3_1517448501_3118;
   wire v3_1517448501_3119;
   wire v3_1517448501_3120;
   wire v3_1517448501_3121;
   wire v3_1517448501_3122;
   wire v3_1517448501_3123;
   wire v3_1517448501_3124;
   wire v3_1517448501_3125;
   wire v3_1517448501_3126;
   wire v3_1517448501_3127;
   wire v3_1517448501_3128;
   wire v3_1517448501_3129;
   wire v3_1517448501_3130;
   wire v3_1517448501_3131;
   wire v3_1517448501_3132;
   wire v3_1517448501_3133;
   wire v3_1517448501_3134;
   wire v3_1517448501_3135;
   wire v3_1517448501_3136;
   wire v3_1517448501_3137;
   wire v3_1517448501_3138;
   wire v3_1517448501_3139;
   wire v3_1517448501_3140;
   wire v3_1517448501_3141;
   wire v3_1517448501_3142;
   wire v3_1517448501_3143;
   wire v3_1517448501_3144;
   wire v3_1517448501_3145;
   wire v3_1517448501_3146;
   wire v3_1517448501_3147;
   wire v3_1517448501_3148;

   // Output Net Declarations
   wire id78;

   // Combinational Assignments
   assign id0 = 1'b0; 
   assign v3_1517448501_70 = 32'b00000000_00000000_00000000_00000111; 
   assign v3_1517448501_71 = 16'b00000000_00000000; 
   assign v3_1517448501_72 = {v_party_responder_0, v3_1517448501_71};
   assign v3_1517448501_73 = 5'b10000; 
   assign v3_1517448501_74 = v3_1517448501_77 ? ~v3_1517448501_76 : v3_1517448501_75;
   assign v3_1517448501_75 = v3_1517448501_72 >> v3_1517448501_73;
   assign v3_1517448501_76 = ~v3_1517448501_72 >> v3_1517448501_73;
   assign v3_1517448501_77 = v3_1517448501_72[31];
   assign v3_1517448501_78 = v3_1517448501_70 == v3_1517448501_74;
   assign v3_1517448501_79 = a_finished_responder_0 & v3_1517448501_78;
   assign v3_1517448501_80 = ~dve_invalid & v3_1517448501_79;
   assign v3_1517448501_82 = 16'b00000110_11101011; 
   assign v3_1517448501_84 = 16'b00000110_01100100; 
   assign v3_1517448501_86 = 16'b00000110_00110111; 
   assign v3_1517448501_88 = 32'b00000000_00000000_00000000_01011010; 
   assign v3_1517448501_89 = {v_party_nonce_responder_2, v3_1517448501_71};
   assign v3_1517448501_90 = v3_1517448501_93 ? ~v3_1517448501_92 : v3_1517448501_91;
   assign v3_1517448501_91 = v3_1517448501_89 >> v3_1517448501_73;
   assign v3_1517448501_92 = ~v3_1517448501_89 >> v3_1517448501_73;
   assign v3_1517448501_93 = v3_1517448501_89[31];
   assign v3_1517448501_94 = v3_1517448501_88 + v3_1517448501_90;
   assign v3_1517448501_95 = 32'b00000000_00000000_00000000_00001111; 
   assign v3_1517448501_96 = {v_party_responder_2, v3_1517448501_71};
   assign v3_1517448501_97 = v3_1517448501_100 ? ~v3_1517448501_99 : v3_1517448501_98;
   assign v3_1517448501_98 = v3_1517448501_96 >> v3_1517448501_73;
   assign v3_1517448501_99 = ~v3_1517448501_96 >> v3_1517448501_73;
   assign v3_1517448501_100 = v3_1517448501_96[31];
   assign v3_1517448501_101 = v3_1517448501_95 * v3_1517448501_97;
   assign v3_1517448501_102 = v3_1517448501_95 * v3_1517448501_101;
   assign v3_1517448501_103 = v3_1517448501_94 + v3_1517448501_102;
   assign v3_1517448501_104 = v3_1517448501_103[15:0];
   assign v3_1517448501_106 = 32'b00000000_00000000_00000000_01001011; 
   assign v3_1517448501_107 = {v_party_nonce_responder_1, v3_1517448501_71};
   assign v3_1517448501_108 = v3_1517448501_111 ? ~v3_1517448501_110 : v3_1517448501_109;
   assign v3_1517448501_109 = v3_1517448501_107 >> v3_1517448501_73;
   assign v3_1517448501_110 = ~v3_1517448501_107 >> v3_1517448501_73;
   assign v3_1517448501_111 = v3_1517448501_107[31];
   assign v3_1517448501_112 = v3_1517448501_106 + v3_1517448501_108;
   assign v3_1517448501_113 = {v_party_responder_1, v3_1517448501_71};
   assign v3_1517448501_114 = v3_1517448501_117 ? ~v3_1517448501_116 : v3_1517448501_115;
   assign v3_1517448501_115 = v3_1517448501_113 >> v3_1517448501_73;
   assign v3_1517448501_116 = ~v3_1517448501_113 >> v3_1517448501_73;
   assign v3_1517448501_117 = v3_1517448501_113[31];
   assign v3_1517448501_118 = v3_1517448501_95 * v3_1517448501_114;
   assign v3_1517448501_119 = v3_1517448501_95 * v3_1517448501_118;
   assign v3_1517448501_120 = v3_1517448501_112 + v3_1517448501_119;
   assign v3_1517448501_121 = v3_1517448501_120[15:0];
   assign v3_1517448501_123 = 32'b00000000_00000000_00000000_00111100; 
   assign v3_1517448501_124 = {v_party_nonce_responder_0, v3_1517448501_71};
   assign v3_1517448501_125 = v3_1517448501_128 ? ~v3_1517448501_127 : v3_1517448501_126;
   assign v3_1517448501_126 = v3_1517448501_124 >> v3_1517448501_73;
   assign v3_1517448501_127 = ~v3_1517448501_124 >> v3_1517448501_73;
   assign v3_1517448501_128 = v3_1517448501_124[31];
   assign v3_1517448501_129 = v3_1517448501_123 + v3_1517448501_125;
   assign v3_1517448501_130 = v3_1517448501_95 * v3_1517448501_74;
   assign v3_1517448501_131 = v3_1517448501_95 * v3_1517448501_130;
   assign v3_1517448501_132 = v3_1517448501_129 + v3_1517448501_131;
   assign v3_1517448501_133 = v3_1517448501_132[15:0];
   assign v3_1517448501_134 = f111 ? v3_1517448501_133 : v_m_initiator_0;
   assign v3_1517448501_135 = f115 ? v3_1517448501_121 : v3_1517448501_134;
   assign v3_1517448501_136 = f119 ? v3_1517448501_104 : v3_1517448501_135;
   assign v3_1517448501_137 = f123 ? v3_1517448501_86 : v3_1517448501_136;
   assign v3_1517448501_138 = f126 ? v3_1517448501_84 : v3_1517448501_137;
   assign v3_1517448501_139 = f129 ? v3_1517448501_82 : v3_1517448501_138;
   assign v3_1517448501_140 = 16'b00000000_00000000; 
   assign v3_1517448501_142 = {v_m_initiator_0, v3_1517448501_71};
   assign v3_1517448501_143 = v3_1517448501_146 ? ~v3_1517448501_145 : v3_1517448501_144;
   assign v3_1517448501_144 = v3_1517448501_142 >> v3_1517448501_73;
   assign v3_1517448501_145 = ~v3_1517448501_142 >> v3_1517448501_73;
   assign v3_1517448501_146 = v3_1517448501_142[31];
   assign v3_1517448501_147 = 32'b00000000_00000000_00000000_11100001; 
   assign v3_1517448501_148 = v3_1517448501_149 ? v3_1517448501_157 : v3_1517448501_156;
   assign v3_1517448501_149 = v3_1517448501_143[31];
   assign v3_1517448501_150 = v3_1517448501_147[31];
   assign v3_1517448501_151 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_152 = ~v3_1517448501_143 + v3_1517448501_151;
   assign v3_1517448501_153 = ~v3_1517448501_147 + v3_1517448501_151;
   assign v3_1517448501_154 = v3_1517448501_149 ? v3_1517448501_152 : v3_1517448501_143;
   assign v3_1517448501_155 = v3_1517448501_150 ? v3_1517448501_153 : v3_1517448501_147;
   assign v3_1517448501_156 = v3_1517448501_154 % v3_1517448501_155;
   assign v3_1517448501_157 = ~v3_1517448501_156 + v3_1517448501_151;
   assign v3_1517448501_158 = v3_1517448501_161 ? v3_1517448501_168 : v3_1517448501_167;
   assign v3_1517448501_159 = v3_1517448501_148[31];
   assign v3_1517448501_160 = v3_1517448501_95[31];
   assign v3_1517448501_161 = v3_1517448501_159 ^ v3_1517448501_160;
   assign v3_1517448501_162 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_163 = ~v3_1517448501_148 + v3_1517448501_162;
   assign v3_1517448501_164 = ~v3_1517448501_95 + v3_1517448501_162;
   assign v3_1517448501_165 = v3_1517448501_159 ? v3_1517448501_163 : v3_1517448501_148;
   assign v3_1517448501_166 = v3_1517448501_160 ? v3_1517448501_164 : v3_1517448501_95;
   assign v3_1517448501_167 = v3_1517448501_165 / v3_1517448501_166;
   assign v3_1517448501_168 = ~v3_1517448501_167 + v3_1517448501_162;
   assign v3_1517448501_169 = v3_1517448501_158[15:0];
   assign v3_1517448501_170 = f000 ? v3_1517448501_169 : v_party_nonce_initiator_0;
   assign v3_1517448501_171 = 16'b00000000_00000000; 
   assign v3_1517448501_178 = f112 ? v3_1517448501_133 : v_m_initiator_1;
   assign v3_1517448501_179 = f116 ? v3_1517448501_121 : v3_1517448501_178;
   assign v3_1517448501_180 = f120 ? v3_1517448501_104 : v3_1517448501_179;
   assign v3_1517448501_181 = f124 ? v3_1517448501_86 : v3_1517448501_180;
   assign v3_1517448501_182 = f127 ? v3_1517448501_84 : v3_1517448501_181;
   assign v3_1517448501_183 = f130 ? v3_1517448501_82 : v3_1517448501_182;
   assign v3_1517448501_184 = 16'b00000000_00000000; 
   assign v3_1517448501_186 = {v_m_initiator_1, v3_1517448501_71};
   assign v3_1517448501_187 = v3_1517448501_190 ? ~v3_1517448501_189 : v3_1517448501_188;
   assign v3_1517448501_188 = v3_1517448501_186 >> v3_1517448501_73;
   assign v3_1517448501_189 = ~v3_1517448501_186 >> v3_1517448501_73;
   assign v3_1517448501_190 = v3_1517448501_186[31];
   assign v3_1517448501_191 = v3_1517448501_192 ? v3_1517448501_200 : v3_1517448501_199;
   assign v3_1517448501_192 = v3_1517448501_187[31];
   assign v3_1517448501_193 = v3_1517448501_147[31];
   assign v3_1517448501_194 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_195 = ~v3_1517448501_187 + v3_1517448501_194;
   assign v3_1517448501_196 = ~v3_1517448501_147 + v3_1517448501_194;
   assign v3_1517448501_197 = v3_1517448501_192 ? v3_1517448501_195 : v3_1517448501_187;
   assign v3_1517448501_198 = v3_1517448501_193 ? v3_1517448501_196 : v3_1517448501_147;
   assign v3_1517448501_199 = v3_1517448501_197 % v3_1517448501_198;
   assign v3_1517448501_200 = ~v3_1517448501_199 + v3_1517448501_194;
   assign v3_1517448501_201 = v3_1517448501_204 ? v3_1517448501_211 : v3_1517448501_210;
   assign v3_1517448501_202 = v3_1517448501_191[31];
   assign v3_1517448501_203 = v3_1517448501_95[31];
   assign v3_1517448501_204 = v3_1517448501_202 ^ v3_1517448501_203;
   assign v3_1517448501_205 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_206 = ~v3_1517448501_191 + v3_1517448501_205;
   assign v3_1517448501_207 = ~v3_1517448501_95 + v3_1517448501_205;
   assign v3_1517448501_208 = v3_1517448501_202 ? v3_1517448501_206 : v3_1517448501_191;
   assign v3_1517448501_209 = v3_1517448501_203 ? v3_1517448501_207 : v3_1517448501_95;
   assign v3_1517448501_210 = v3_1517448501_208 / v3_1517448501_209;
   assign v3_1517448501_211 = ~v3_1517448501_210 + v3_1517448501_205;
   assign v3_1517448501_212 = v3_1517448501_201[15:0];
   assign v3_1517448501_213 = f002 ? v3_1517448501_212 : v_party_nonce_initiator_1;
   assign v3_1517448501_214 = 16'b00000000_00000000; 
   assign v3_1517448501_221 = f113 ? v3_1517448501_133 : v_m_initiator_2;
   assign v3_1517448501_222 = f117 ? v3_1517448501_121 : v3_1517448501_221;
   assign v3_1517448501_223 = f121 ? v3_1517448501_104 : v3_1517448501_222;
   assign v3_1517448501_224 = f125 ? v3_1517448501_86 : v3_1517448501_223;
   assign v3_1517448501_225 = f128 ? v3_1517448501_84 : v3_1517448501_224;
   assign v3_1517448501_226 = f131 ? v3_1517448501_82 : v3_1517448501_225;
   assign v3_1517448501_227 = 16'b00000000_00000000; 
   assign v3_1517448501_229 = {v_m_initiator_2, v3_1517448501_71};
   assign v3_1517448501_230 = v3_1517448501_233 ? ~v3_1517448501_232 : v3_1517448501_231;
   assign v3_1517448501_231 = v3_1517448501_229 >> v3_1517448501_73;
   assign v3_1517448501_232 = ~v3_1517448501_229 >> v3_1517448501_73;
   assign v3_1517448501_233 = v3_1517448501_229[31];
   assign v3_1517448501_234 = v3_1517448501_235 ? v3_1517448501_243 : v3_1517448501_242;
   assign v3_1517448501_235 = v3_1517448501_230[31];
   assign v3_1517448501_236 = v3_1517448501_147[31];
   assign v3_1517448501_237 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_238 = ~v3_1517448501_230 + v3_1517448501_237;
   assign v3_1517448501_239 = ~v3_1517448501_147 + v3_1517448501_237;
   assign v3_1517448501_240 = v3_1517448501_235 ? v3_1517448501_238 : v3_1517448501_230;
   assign v3_1517448501_241 = v3_1517448501_236 ? v3_1517448501_239 : v3_1517448501_147;
   assign v3_1517448501_242 = v3_1517448501_240 % v3_1517448501_241;
   assign v3_1517448501_243 = ~v3_1517448501_242 + v3_1517448501_237;
   assign v3_1517448501_244 = v3_1517448501_247 ? v3_1517448501_254 : v3_1517448501_253;
   assign v3_1517448501_245 = v3_1517448501_234[31];
   assign v3_1517448501_246 = v3_1517448501_95[31];
   assign v3_1517448501_247 = v3_1517448501_245 ^ v3_1517448501_246;
   assign v3_1517448501_248 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_249 = ~v3_1517448501_234 + v3_1517448501_248;
   assign v3_1517448501_250 = ~v3_1517448501_95 + v3_1517448501_248;
   assign v3_1517448501_251 = v3_1517448501_245 ? v3_1517448501_249 : v3_1517448501_234;
   assign v3_1517448501_252 = v3_1517448501_246 ? v3_1517448501_250 : v3_1517448501_95;
   assign v3_1517448501_253 = v3_1517448501_251 / v3_1517448501_252;
   assign v3_1517448501_254 = ~v3_1517448501_253 + v3_1517448501_248;
   assign v3_1517448501_255 = v3_1517448501_244[15:0];
   assign v3_1517448501_256 = f004 ? v3_1517448501_255 : v_party_nonce_initiator_2;
   assign v3_1517448501_257 = 16'b00000000_00000000; 
   assign v3_1517448501_259 = 16'b00000000_10011010; 
   assign v3_1517448501_261 = 32'b00000000_00000000_00000000_10110100; 
   assign v3_1517448501_262 = {v_party_nonce_initiator_2, v3_1517448501_71};
   assign v3_1517448501_263 = v3_1517448501_266 ? ~v3_1517448501_265 : v3_1517448501_264;
   assign v3_1517448501_264 = v3_1517448501_262 >> v3_1517448501_73;
   assign v3_1517448501_265 = ~v3_1517448501_262 >> v3_1517448501_73;
   assign v3_1517448501_266 = v3_1517448501_262[31];
   assign v3_1517448501_267 = v3_1517448501_261 + v3_1517448501_263;
   assign v3_1517448501_268 = v3_1517448501_267[15:0];
   assign v3_1517448501_270 = 32'b00000000_00000000_00000000_10100101; 
   assign v3_1517448501_271 = {v_party_nonce_initiator_1, v3_1517448501_71};
   assign v3_1517448501_272 = v3_1517448501_275 ? ~v3_1517448501_274 : v3_1517448501_273;
   assign v3_1517448501_273 = v3_1517448501_271 >> v3_1517448501_73;
   assign v3_1517448501_274 = ~v3_1517448501_271 >> v3_1517448501_73;
   assign v3_1517448501_275 = v3_1517448501_271[31];
   assign v3_1517448501_276 = v3_1517448501_270 + v3_1517448501_272;
   assign v3_1517448501_277 = v3_1517448501_276[15:0];
   assign v3_1517448501_279 = 32'b00000000_00000000_00000000_10010110; 
   assign v3_1517448501_280 = {v_party_nonce_initiator_0, v3_1517448501_71};
   assign v3_1517448501_281 = v3_1517448501_284 ? ~v3_1517448501_283 : v3_1517448501_282;
   assign v3_1517448501_282 = v3_1517448501_280 >> v3_1517448501_73;
   assign v3_1517448501_283 = ~v3_1517448501_280 >> v3_1517448501_73;
   assign v3_1517448501_284 = v3_1517448501_280[31];
   assign v3_1517448501_285 = v3_1517448501_279 + v3_1517448501_281;
   assign v3_1517448501_286 = v3_1517448501_285[15:0];
   assign v3_1517448501_288 = 16'b00001000_11111011; 
   assign v3_1517448501_290 = 16'b00001001_01100100; 
   assign v3_1517448501_292 = 16'b00001001_00110111; 
   assign v3_1517448501_294 = 16'b00001000_11111000; 
   assign v3_1517448501_296 = 16'b00001001_01100001; 
   assign v3_1517448501_298 = 16'b00001001_00110100; 
   assign v3_1517448501_300 = 16'b00000110_01010101; 
   assign v3_1517448501_302 = 16'b00000110_10111110; 
   assign v3_1517448501_304 = 16'b00000110_10010001; 
   assign v3_1517448501_306 = 16'b00001000_11111010; 
   assign v3_1517448501_308 = 16'b00001001_01100011; 
   assign v3_1517448501_310 = 16'b00001001_00110110; 
   assign v3_1517448501_312 = 16'b00001001_00000001; 
   assign v3_1517448501_314 = 16'b00001001_01101010; 
   assign v3_1517448501_316 = 16'b00001001_00111101; 
   assign v3_1517448501_318 = 16'b00001000_11111110; 
   assign v3_1517448501_320 = 16'b00001001_01100111; 
   assign v3_1517448501_322 = 16'b00001001_00111010; 
   assign v3_1517448501_324 = 16'b00001001_00000100; 
   assign v3_1517448501_326 = 16'b00001001_01101101; 
   assign v3_1517448501_328 = 16'b00001001_01000000; 
   assign v3_1517448501_330 = 16'b00001011_00010110; 
   assign v3_1517448501_332 = 16'b00001010_00100101; 
   assign v3_1517448501_334 = f036 ? v3_1517448501_298 : v_m_responder_0;
   assign v3_1517448501_335 = f040 ? v3_1517448501_332 : v3_1517448501_334;
   assign v3_1517448501_336 = f044 ? v3_1517448501_330 : v3_1517448501_335;
   assign v3_1517448501_337 = f048 ? v3_1517448501_328 : v3_1517448501_336;
   assign v3_1517448501_338 = f051 ? v3_1517448501_326 : v3_1517448501_337;
   assign v3_1517448501_339 = f054 ? v3_1517448501_324 : v3_1517448501_338;
   assign v3_1517448501_340 = f057 ? v3_1517448501_322 : v3_1517448501_339;
   assign v3_1517448501_341 = f060 ? v3_1517448501_320 : v3_1517448501_340;
   assign v3_1517448501_342 = f063 ? v3_1517448501_318 : v3_1517448501_341;
   assign v3_1517448501_343 = f066 ? v3_1517448501_316 : v3_1517448501_342;
   assign v3_1517448501_344 = f069 ? v3_1517448501_314 : v3_1517448501_343;
   assign v3_1517448501_345 = f072 ? v3_1517448501_312 : v3_1517448501_344;
   assign v3_1517448501_346 = f075 ? v3_1517448501_310 : v3_1517448501_345;
   assign v3_1517448501_347 = f078 ? v3_1517448501_308 : v3_1517448501_346;
   assign v3_1517448501_348 = f081 ? v3_1517448501_306 : v3_1517448501_347;
   assign v3_1517448501_349 = f084 ? v3_1517448501_304 : v3_1517448501_348;
   assign v3_1517448501_350 = f087 ? v3_1517448501_302 : v3_1517448501_349;
   assign v3_1517448501_351 = f090 ? v3_1517448501_300 : v3_1517448501_350;
   assign v3_1517448501_352 = f093 ? v3_1517448501_298 : v3_1517448501_351;
   assign v3_1517448501_353 = f096 ? v3_1517448501_296 : v3_1517448501_352;
   assign v3_1517448501_354 = f099 ? v3_1517448501_294 : v3_1517448501_353;
   assign v3_1517448501_355 = f102 ? v3_1517448501_292 : v3_1517448501_354;
   assign v3_1517448501_356 = f105 ? v3_1517448501_290 : v3_1517448501_355;
   assign v3_1517448501_357 = f108 ? v3_1517448501_288 : v3_1517448501_356;
   assign v3_1517448501_358 = f132 ? v3_1517448501_286 : v3_1517448501_357;
   assign v3_1517448501_359 = f136 ? v3_1517448501_277 : v3_1517448501_358;
   assign v3_1517448501_360 = f140 ? v3_1517448501_268 : v3_1517448501_359;
   assign v3_1517448501_361 = f144 ? v3_1517448501_259 : v3_1517448501_360;
   assign v3_1517448501_362 = 16'b00000000_00000000; 
   assign v3_1517448501_364 = {v_m_responder_0, v3_1517448501_71};
   assign v3_1517448501_365 = v3_1517448501_368 ? ~v3_1517448501_367 : v3_1517448501_366;
   assign v3_1517448501_366 = v3_1517448501_364 >> v3_1517448501_73;
   assign v3_1517448501_367 = ~v3_1517448501_364 >> v3_1517448501_73;
   assign v3_1517448501_368 = v3_1517448501_364[31];
   assign v3_1517448501_369 = v3_1517448501_370 ? v3_1517448501_378 : v3_1517448501_377;
   assign v3_1517448501_370 = v3_1517448501_365[31];
   assign v3_1517448501_371 = v3_1517448501_147[31];
   assign v3_1517448501_372 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_373 = ~v3_1517448501_365 + v3_1517448501_372;
   assign v3_1517448501_374 = ~v3_1517448501_147 + v3_1517448501_372;
   assign v3_1517448501_375 = v3_1517448501_370 ? v3_1517448501_373 : v3_1517448501_365;
   assign v3_1517448501_376 = v3_1517448501_371 ? v3_1517448501_374 : v3_1517448501_147;
   assign v3_1517448501_377 = v3_1517448501_375 % v3_1517448501_376;
   assign v3_1517448501_378 = ~v3_1517448501_377 + v3_1517448501_372;
   assign v3_1517448501_379 = v3_1517448501_382 ? v3_1517448501_389 : v3_1517448501_388;
   assign v3_1517448501_380 = v3_1517448501_369[31];
   assign v3_1517448501_381 = v3_1517448501_95[31];
   assign v3_1517448501_382 = v3_1517448501_380 ^ v3_1517448501_381;
   assign v3_1517448501_383 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_384 = ~v3_1517448501_369 + v3_1517448501_383;
   assign v3_1517448501_385 = ~v3_1517448501_95 + v3_1517448501_383;
   assign v3_1517448501_386 = v3_1517448501_380 ? v3_1517448501_384 : v3_1517448501_369;
   assign v3_1517448501_387 = v3_1517448501_381 ? v3_1517448501_385 : v3_1517448501_95;
   assign v3_1517448501_388 = v3_1517448501_386 / v3_1517448501_387;
   assign v3_1517448501_389 = ~v3_1517448501_388 + v3_1517448501_383;
   assign v3_1517448501_390 = v3_1517448501_379[15:0];
   assign v3_1517448501_391 = f006 ? v3_1517448501_390 : v_party_responder_0;
   assign v3_1517448501_392 = 16'b00000000_00000000; 
   assign v3_1517448501_393 = v3_1517448501_394 ? v3_1517448501_402 : v3_1517448501_401;
   assign v3_1517448501_394 = v3_1517448501_365[31];
   assign v3_1517448501_395 = v3_1517448501_95[31];
   assign v3_1517448501_396 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_397 = ~v3_1517448501_365 + v3_1517448501_396;
   assign v3_1517448501_398 = ~v3_1517448501_95 + v3_1517448501_396;
   assign v3_1517448501_399 = v3_1517448501_394 ? v3_1517448501_397 : v3_1517448501_365;
   assign v3_1517448501_400 = v3_1517448501_395 ? v3_1517448501_398 : v3_1517448501_95;
   assign v3_1517448501_401 = v3_1517448501_399 % v3_1517448501_400;
   assign v3_1517448501_402 = ~v3_1517448501_401 + v3_1517448501_396;
   assign v3_1517448501_403 = v3_1517448501_393[15:0];
   assign v3_1517448501_404 = f006 ? v3_1517448501_403 : v_party_nonce_responder_0;
   assign v3_1517448501_405 = 16'b00000000_00000000; 
   assign v3_1517448501_434 = f037 ? v3_1517448501_298 : v_m_responder_1;
   assign v3_1517448501_435 = f041 ? v3_1517448501_332 : v3_1517448501_434;
   assign v3_1517448501_436 = f045 ? v3_1517448501_330 : v3_1517448501_435;
   assign v3_1517448501_437 = f049 ? v3_1517448501_328 : v3_1517448501_436;
   assign v3_1517448501_438 = f052 ? v3_1517448501_326 : v3_1517448501_437;
   assign v3_1517448501_439 = f055 ? v3_1517448501_324 : v3_1517448501_438;
   assign v3_1517448501_440 = f058 ? v3_1517448501_322 : v3_1517448501_439;
   assign v3_1517448501_441 = f061 ? v3_1517448501_320 : v3_1517448501_440;
   assign v3_1517448501_442 = f064 ? v3_1517448501_318 : v3_1517448501_441;
   assign v3_1517448501_443 = f067 ? v3_1517448501_316 : v3_1517448501_442;
   assign v3_1517448501_444 = f070 ? v3_1517448501_314 : v3_1517448501_443;
   assign v3_1517448501_445 = f073 ? v3_1517448501_312 : v3_1517448501_444;
   assign v3_1517448501_446 = f076 ? v3_1517448501_310 : v3_1517448501_445;
   assign v3_1517448501_447 = f079 ? v3_1517448501_308 : v3_1517448501_446;
   assign v3_1517448501_448 = f082 ? v3_1517448501_306 : v3_1517448501_447;
   assign v3_1517448501_449 = f085 ? v3_1517448501_304 : v3_1517448501_448;
   assign v3_1517448501_450 = f088 ? v3_1517448501_302 : v3_1517448501_449;
   assign v3_1517448501_451 = f091 ? v3_1517448501_300 : v3_1517448501_450;
   assign v3_1517448501_452 = f094 ? v3_1517448501_298 : v3_1517448501_451;
   assign v3_1517448501_453 = f097 ? v3_1517448501_296 : v3_1517448501_452;
   assign v3_1517448501_454 = f100 ? v3_1517448501_294 : v3_1517448501_453;
   assign v3_1517448501_455 = f103 ? v3_1517448501_292 : v3_1517448501_454;
   assign v3_1517448501_456 = f106 ? v3_1517448501_290 : v3_1517448501_455;
   assign v3_1517448501_457 = f109 ? v3_1517448501_288 : v3_1517448501_456;
   assign v3_1517448501_458 = f133 ? v3_1517448501_286 : v3_1517448501_457;
   assign v3_1517448501_459 = f137 ? v3_1517448501_277 : v3_1517448501_458;
   assign v3_1517448501_460 = f141 ? v3_1517448501_268 : v3_1517448501_459;
   assign v3_1517448501_461 = f145 ? v3_1517448501_259 : v3_1517448501_460;
   assign v3_1517448501_462 = 16'b00000000_00000000; 
   assign v3_1517448501_464 = {v_m_responder_1, v3_1517448501_71};
   assign v3_1517448501_465 = v3_1517448501_468 ? ~v3_1517448501_467 : v3_1517448501_466;
   assign v3_1517448501_466 = v3_1517448501_464 >> v3_1517448501_73;
   assign v3_1517448501_467 = ~v3_1517448501_464 >> v3_1517448501_73;
   assign v3_1517448501_468 = v3_1517448501_464[31];
   assign v3_1517448501_469 = v3_1517448501_470 ? v3_1517448501_478 : v3_1517448501_477;
   assign v3_1517448501_470 = v3_1517448501_465[31];
   assign v3_1517448501_471 = v3_1517448501_147[31];
   assign v3_1517448501_472 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_473 = ~v3_1517448501_465 + v3_1517448501_472;
   assign v3_1517448501_474 = ~v3_1517448501_147 + v3_1517448501_472;
   assign v3_1517448501_475 = v3_1517448501_470 ? v3_1517448501_473 : v3_1517448501_465;
   assign v3_1517448501_476 = v3_1517448501_471 ? v3_1517448501_474 : v3_1517448501_147;
   assign v3_1517448501_477 = v3_1517448501_475 % v3_1517448501_476;
   assign v3_1517448501_478 = ~v3_1517448501_477 + v3_1517448501_472;
   assign v3_1517448501_479 = v3_1517448501_482 ? v3_1517448501_489 : v3_1517448501_488;
   assign v3_1517448501_480 = v3_1517448501_469[31];
   assign v3_1517448501_481 = v3_1517448501_95[31];
   assign v3_1517448501_482 = v3_1517448501_480 ^ v3_1517448501_481;
   assign v3_1517448501_483 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_484 = ~v3_1517448501_469 + v3_1517448501_483;
   assign v3_1517448501_485 = ~v3_1517448501_95 + v3_1517448501_483;
   assign v3_1517448501_486 = v3_1517448501_480 ? v3_1517448501_484 : v3_1517448501_469;
   assign v3_1517448501_487 = v3_1517448501_481 ? v3_1517448501_485 : v3_1517448501_95;
   assign v3_1517448501_488 = v3_1517448501_486 / v3_1517448501_487;
   assign v3_1517448501_489 = ~v3_1517448501_488 + v3_1517448501_483;
   assign v3_1517448501_490 = v3_1517448501_479[15:0];
   assign v3_1517448501_491 = f010 ? v3_1517448501_490 : v_party_responder_1;
   assign v3_1517448501_492 = 16'b00000000_00000000; 
   assign v3_1517448501_493 = v3_1517448501_494 ? v3_1517448501_502 : v3_1517448501_501;
   assign v3_1517448501_494 = v3_1517448501_465[31];
   assign v3_1517448501_495 = v3_1517448501_95[31];
   assign v3_1517448501_496 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_497 = ~v3_1517448501_465 + v3_1517448501_496;
   assign v3_1517448501_498 = ~v3_1517448501_95 + v3_1517448501_496;
   assign v3_1517448501_499 = v3_1517448501_494 ? v3_1517448501_497 : v3_1517448501_465;
   assign v3_1517448501_500 = v3_1517448501_495 ? v3_1517448501_498 : v3_1517448501_95;
   assign v3_1517448501_501 = v3_1517448501_499 % v3_1517448501_500;
   assign v3_1517448501_502 = ~v3_1517448501_501 + v3_1517448501_496;
   assign v3_1517448501_503 = v3_1517448501_493[15:0];
   assign v3_1517448501_504 = f010 ? v3_1517448501_503 : v_party_nonce_responder_1;
   assign v3_1517448501_505 = 16'b00000000_00000000; 
   assign v3_1517448501_534 = f038 ? v3_1517448501_298 : v_m_responder_2;
   assign v3_1517448501_535 = f042 ? v3_1517448501_332 : v3_1517448501_534;
   assign v3_1517448501_536 = f046 ? v3_1517448501_330 : v3_1517448501_535;
   assign v3_1517448501_537 = f050 ? v3_1517448501_328 : v3_1517448501_536;
   assign v3_1517448501_538 = f053 ? v3_1517448501_326 : v3_1517448501_537;
   assign v3_1517448501_539 = f056 ? v3_1517448501_324 : v3_1517448501_538;
   assign v3_1517448501_540 = f059 ? v3_1517448501_322 : v3_1517448501_539;
   assign v3_1517448501_541 = f062 ? v3_1517448501_320 : v3_1517448501_540;
   assign v3_1517448501_542 = f065 ? v3_1517448501_318 : v3_1517448501_541;
   assign v3_1517448501_543 = f068 ? v3_1517448501_316 : v3_1517448501_542;
   assign v3_1517448501_544 = f071 ? v3_1517448501_314 : v3_1517448501_543;
   assign v3_1517448501_545 = f074 ? v3_1517448501_312 : v3_1517448501_544;
   assign v3_1517448501_546 = f077 ? v3_1517448501_310 : v3_1517448501_545;
   assign v3_1517448501_547 = f080 ? v3_1517448501_308 : v3_1517448501_546;
   assign v3_1517448501_548 = f083 ? v3_1517448501_306 : v3_1517448501_547;
   assign v3_1517448501_549 = f086 ? v3_1517448501_304 : v3_1517448501_548;
   assign v3_1517448501_550 = f089 ? v3_1517448501_302 : v3_1517448501_549;
   assign v3_1517448501_551 = f092 ? v3_1517448501_300 : v3_1517448501_550;
   assign v3_1517448501_552 = f095 ? v3_1517448501_298 : v3_1517448501_551;
   assign v3_1517448501_553 = f098 ? v3_1517448501_296 : v3_1517448501_552;
   assign v3_1517448501_554 = f101 ? v3_1517448501_294 : v3_1517448501_553;
   assign v3_1517448501_555 = f104 ? v3_1517448501_292 : v3_1517448501_554;
   assign v3_1517448501_556 = f107 ? v3_1517448501_290 : v3_1517448501_555;
   assign v3_1517448501_557 = f110 ? v3_1517448501_288 : v3_1517448501_556;
   assign v3_1517448501_558 = f134 ? v3_1517448501_286 : v3_1517448501_557;
   assign v3_1517448501_559 = f138 ? v3_1517448501_277 : v3_1517448501_558;
   assign v3_1517448501_560 = f142 ? v3_1517448501_268 : v3_1517448501_559;
   assign v3_1517448501_561 = f146 ? v3_1517448501_259 : v3_1517448501_560;
   assign v3_1517448501_562 = 16'b00000000_00000000; 
   assign v3_1517448501_564 = {v_m_responder_2, v3_1517448501_71};
   assign v3_1517448501_565 = v3_1517448501_568 ? ~v3_1517448501_567 : v3_1517448501_566;
   assign v3_1517448501_566 = v3_1517448501_564 >> v3_1517448501_73;
   assign v3_1517448501_567 = ~v3_1517448501_564 >> v3_1517448501_73;
   assign v3_1517448501_568 = v3_1517448501_564[31];
   assign v3_1517448501_569 = v3_1517448501_570 ? v3_1517448501_578 : v3_1517448501_577;
   assign v3_1517448501_570 = v3_1517448501_565[31];
   assign v3_1517448501_571 = v3_1517448501_147[31];
   assign v3_1517448501_572 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_573 = ~v3_1517448501_565 + v3_1517448501_572;
   assign v3_1517448501_574 = ~v3_1517448501_147 + v3_1517448501_572;
   assign v3_1517448501_575 = v3_1517448501_570 ? v3_1517448501_573 : v3_1517448501_565;
   assign v3_1517448501_576 = v3_1517448501_571 ? v3_1517448501_574 : v3_1517448501_147;
   assign v3_1517448501_577 = v3_1517448501_575 % v3_1517448501_576;
   assign v3_1517448501_578 = ~v3_1517448501_577 + v3_1517448501_572;
   assign v3_1517448501_579 = v3_1517448501_582 ? v3_1517448501_589 : v3_1517448501_588;
   assign v3_1517448501_580 = v3_1517448501_569[31];
   assign v3_1517448501_581 = v3_1517448501_95[31];
   assign v3_1517448501_582 = v3_1517448501_580 ^ v3_1517448501_581;
   assign v3_1517448501_583 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_584 = ~v3_1517448501_569 + v3_1517448501_583;
   assign v3_1517448501_585 = ~v3_1517448501_95 + v3_1517448501_583;
   assign v3_1517448501_586 = v3_1517448501_580 ? v3_1517448501_584 : v3_1517448501_569;
   assign v3_1517448501_587 = v3_1517448501_581 ? v3_1517448501_585 : v3_1517448501_95;
   assign v3_1517448501_588 = v3_1517448501_586 / v3_1517448501_587;
   assign v3_1517448501_589 = ~v3_1517448501_588 + v3_1517448501_583;
   assign v3_1517448501_590 = v3_1517448501_579[15:0];
   assign v3_1517448501_591 = f014 ? v3_1517448501_590 : v_party_responder_2;
   assign v3_1517448501_592 = 16'b00000000_00000000; 
   assign v3_1517448501_593 = v3_1517448501_594 ? v3_1517448501_602 : v3_1517448501_601;
   assign v3_1517448501_594 = v3_1517448501_565[31];
   assign v3_1517448501_595 = v3_1517448501_95[31];
   assign v3_1517448501_596 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_597 = ~v3_1517448501_565 + v3_1517448501_596;
   assign v3_1517448501_598 = ~v3_1517448501_95 + v3_1517448501_596;
   assign v3_1517448501_599 = v3_1517448501_594 ? v3_1517448501_597 : v3_1517448501_565;
   assign v3_1517448501_600 = v3_1517448501_595 ? v3_1517448501_598 : v3_1517448501_95;
   assign v3_1517448501_601 = v3_1517448501_599 % v3_1517448501_600;
   assign v3_1517448501_602 = ~v3_1517448501_601 + v3_1517448501_596;
   assign v3_1517448501_603 = v3_1517448501_593[15:0];
   assign v3_1517448501_604 = f014 ? v3_1517448501_603 : v_party_nonce_responder_2;
   assign v3_1517448501_605 = 16'b00000000_00000000; 
   assign v3_1517448501_607 = 8'b00000001; 
   assign v3_1517448501_609 = f021 ? v3_1517448501_607 : v_kNa;
   assign v3_1517448501_610 = f031 ? v3_1517448501_607 : v3_1517448501_609;
   assign v3_1517448501_611 = 8'b00000000; 
   assign v3_1517448501_614 = f022 ? v3_1517448501_607 : v_kNb;
   assign v3_1517448501_615 = f032 ? v3_1517448501_607 : v3_1517448501_614;
   assign v3_1517448501_616 = 8'b00000000; 
   assign v3_1517448501_618 = f027 ? v3_1517448501_607 : v_k_Na_Nb__A;
   assign v3_1517448501_619 = 8'b00000000; 
   assign v3_1517448501_621 = f026 ? v3_1517448501_607 : v_k_Na_A__B;
   assign v3_1517448501_622 = 8'b00000000; 
   assign v3_1517448501_625 = f024 ? v3_1517448501_607 : v_k_Nb__B;
   assign v3_1517448501_626 = f034 ? v3_1517448501_607 : v3_1517448501_625;
   assign v3_1517448501_627 = 8'b00000000; 
   assign v3_1517448501_637 = f039 ? v3_1517448501_298 : v_m_intruder;
   assign v3_1517448501_638 = f043 ? v3_1517448501_332 : v3_1517448501_637;
   assign v3_1517448501_639 = f047 ? v3_1517448501_330 : v3_1517448501_638;
   assign v3_1517448501_640 = f114 ? v3_1517448501_133 : v3_1517448501_639;
   assign v3_1517448501_641 = f118 ? v3_1517448501_121 : v3_1517448501_640;
   assign v3_1517448501_642 = f122 ? v3_1517448501_104 : v3_1517448501_641;
   assign v3_1517448501_643 = f135 ? v3_1517448501_286 : v3_1517448501_642;
   assign v3_1517448501_644 = f139 ? v3_1517448501_277 : v3_1517448501_643;
   assign v3_1517448501_645 = f143 ? v3_1517448501_268 : v3_1517448501_644;
   assign v3_1517448501_646 = 16'b00000000_00000000; 
   assign v3_1517448501_647 = ~a_start_initiator_0 & ~f036;
   assign v3_1517448501_648 = v3_1517448501_647 & ~f037;
   assign v3_1517448501_649 = v3_1517448501_648 & ~f038;
   assign v3_1517448501_650 = v3_1517448501_649 & ~f039;
   assign v3_1517448501_651 = 1'b0; 
   assign v3_1517448501_652 = ~v3_1517448501_653;
   assign v3_1517448501_653 = ~a_wait_resp_initiator_0 & ~f036;
   assign v3_1517448501_654 = ~v3_1517448501_655;
   assign v3_1517448501_655 = ~v3_1517448501_652 & ~f037;
   assign v3_1517448501_656 = ~v3_1517448501_657;
   assign v3_1517448501_657 = ~v3_1517448501_654 & ~f038;
   assign v3_1517448501_658 = ~v3_1517448501_659;
   assign v3_1517448501_659 = ~v3_1517448501_656 & ~f039;
   assign v3_1517448501_660 = v3_1517448501_658 & ~f111;
   assign v3_1517448501_661 = v3_1517448501_660 & ~f115;
   assign v3_1517448501_662 = v3_1517448501_661 & ~f119;
   assign v3_1517448501_663 = v3_1517448501_662 & ~f123;
   assign v3_1517448501_664 = v3_1517448501_663 & ~f126;
   assign v3_1517448501_665 = v3_1517448501_664 & ~f129;
   assign v3_1517448501_666 = 1'b0; 
   assign v3_1517448501_667 = a_got_resp_initiator_0 & ~f000;
   assign v3_1517448501_669 = v3_1517448501_667 & ~f001;
   assign v3_1517448501_670 = ~v3_1517448501_671;
   assign v3_1517448501_671 = ~v3_1517448501_669 & ~f111;
   assign v3_1517448501_672 = ~v3_1517448501_673;
   assign v3_1517448501_673 = ~v3_1517448501_670 & ~f115;
   assign v3_1517448501_674 = ~v3_1517448501_675;
   assign v3_1517448501_675 = ~v3_1517448501_672 & ~f119;
   assign v3_1517448501_676 = ~v3_1517448501_677;
   assign v3_1517448501_677 = ~v3_1517448501_674 & ~f123;
   assign v3_1517448501_678 = ~v3_1517448501_679;
   assign v3_1517448501_679 = ~v3_1517448501_676 & ~f126;
   assign v3_1517448501_680 = ~v3_1517448501_681;
   assign v3_1517448501_681 = ~v3_1517448501_678 & ~f129;
   assign v3_1517448501_682 = 1'b0; 
   assign v3_1517448501_683 = ~v3_1517448501_684;
   assign v3_1517448501_684 = ~a_commited_initiator_0 & ~f000;
   assign v3_1517448501_685 = v3_1517448501_683 & ~f132;
   assign v3_1517448501_686 = v3_1517448501_685 & ~f133;
   assign v3_1517448501_687 = v3_1517448501_686 & ~f134;
   assign v3_1517448501_688 = v3_1517448501_687 & ~f135;
   assign v3_1517448501_689 = 1'b0; 
   assign v3_1517448501_690 = ~v3_1517448501_691;
   assign v3_1517448501_691 = ~a_finished_initiator_0 & ~f132;
   assign v3_1517448501_692 = ~v3_1517448501_693;
   assign v3_1517448501_693 = ~v3_1517448501_690 & ~f133;
   assign v3_1517448501_694 = ~v3_1517448501_695;
   assign v3_1517448501_695 = ~v3_1517448501_692 & ~f134;
   assign v3_1517448501_696 = ~v3_1517448501_697;
   assign v3_1517448501_697 = ~v3_1517448501_694 & ~f135;
   assign v3_1517448501_698 = 1'b0; 
   assign v3_1517448501_699 = ~v3_1517448501_700;
   assign v3_1517448501_700 = ~a_corrupted_initiator_0 & ~f001;
   assign v3_1517448501_701 = 1'b0; 
   assign v3_1517448501_702 = ~a_start_initiator_1 & ~f040;
   assign v3_1517448501_703 = v3_1517448501_702 & ~f041;
   assign v3_1517448501_704 = v3_1517448501_703 & ~f042;
   assign v3_1517448501_705 = v3_1517448501_704 & ~f043;
   assign v3_1517448501_706 = 1'b0; 
   assign v3_1517448501_707 = ~v3_1517448501_708;
   assign v3_1517448501_708 = ~a_wait_resp_initiator_1 & ~f040;
   assign v3_1517448501_709 = ~v3_1517448501_710;
   assign v3_1517448501_710 = ~v3_1517448501_707 & ~f041;
   assign v3_1517448501_711 = ~v3_1517448501_712;
   assign v3_1517448501_712 = ~v3_1517448501_709 & ~f042;
   assign v3_1517448501_713 = ~v3_1517448501_714;
   assign v3_1517448501_714 = ~v3_1517448501_711 & ~f043;
   assign v3_1517448501_715 = v3_1517448501_713 & ~f112;
   assign v3_1517448501_716 = v3_1517448501_715 & ~f116;
   assign v3_1517448501_717 = v3_1517448501_716 & ~f120;
   assign v3_1517448501_718 = v3_1517448501_717 & ~f124;
   assign v3_1517448501_719 = v3_1517448501_718 & ~f127;
   assign v3_1517448501_720 = v3_1517448501_719 & ~f130;
   assign v3_1517448501_721 = 1'b0; 
   assign v3_1517448501_722 = a_got_resp_initiator_1 & ~f002;
   assign v3_1517448501_724 = v3_1517448501_722 & ~f003;
   assign v3_1517448501_725 = ~v3_1517448501_726;
   assign v3_1517448501_726 = ~v3_1517448501_724 & ~f112;
   assign v3_1517448501_727 = ~v3_1517448501_728;
   assign v3_1517448501_728 = ~v3_1517448501_725 & ~f116;
   assign v3_1517448501_729 = ~v3_1517448501_730;
   assign v3_1517448501_730 = ~v3_1517448501_727 & ~f120;
   assign v3_1517448501_731 = ~v3_1517448501_732;
   assign v3_1517448501_732 = ~v3_1517448501_729 & ~f124;
   assign v3_1517448501_733 = ~v3_1517448501_734;
   assign v3_1517448501_734 = ~v3_1517448501_731 & ~f127;
   assign v3_1517448501_735 = ~v3_1517448501_736;
   assign v3_1517448501_736 = ~v3_1517448501_733 & ~f130;
   assign v3_1517448501_737 = 1'b0; 
   assign v3_1517448501_738 = ~v3_1517448501_739;
   assign v3_1517448501_739 = ~a_commited_initiator_1 & ~f002;
   assign v3_1517448501_740 = v3_1517448501_738 & ~f136;
   assign v3_1517448501_741 = v3_1517448501_740 & ~f137;
   assign v3_1517448501_742 = v3_1517448501_741 & ~f138;
   assign v3_1517448501_743 = v3_1517448501_742 & ~f139;
   assign v3_1517448501_744 = 1'b0; 
   assign v3_1517448501_745 = ~v3_1517448501_746;
   assign v3_1517448501_746 = ~a_finished_initiator_1 & ~f136;
   assign v3_1517448501_747 = ~v3_1517448501_748;
   assign v3_1517448501_748 = ~v3_1517448501_745 & ~f137;
   assign v3_1517448501_749 = ~v3_1517448501_750;
   assign v3_1517448501_750 = ~v3_1517448501_747 & ~f138;
   assign v3_1517448501_751 = ~v3_1517448501_752;
   assign v3_1517448501_752 = ~v3_1517448501_749 & ~f139;
   assign v3_1517448501_753 = 1'b0; 
   assign v3_1517448501_754 = ~v3_1517448501_755;
   assign v3_1517448501_755 = ~a_corrupted_initiator_1 & ~f003;
   assign v3_1517448501_756 = 1'b0; 
   assign v3_1517448501_757 = ~a_start_initiator_2 & ~f044;
   assign v3_1517448501_758 = v3_1517448501_757 & ~f045;
   assign v3_1517448501_759 = v3_1517448501_758 & ~f046;
   assign v3_1517448501_760 = v3_1517448501_759 & ~f047;
   assign v3_1517448501_761 = 1'b0; 
   assign v3_1517448501_762 = ~v3_1517448501_763;
   assign v3_1517448501_763 = ~a_wait_resp_initiator_2 & ~f044;
   assign v3_1517448501_764 = ~v3_1517448501_765;
   assign v3_1517448501_765 = ~v3_1517448501_762 & ~f045;
   assign v3_1517448501_766 = ~v3_1517448501_767;
   assign v3_1517448501_767 = ~v3_1517448501_764 & ~f046;
   assign v3_1517448501_768 = ~v3_1517448501_769;
   assign v3_1517448501_769 = ~v3_1517448501_766 & ~f047;
   assign v3_1517448501_770 = v3_1517448501_768 & ~f113;
   assign v3_1517448501_771 = v3_1517448501_770 & ~f117;
   assign v3_1517448501_772 = v3_1517448501_771 & ~f121;
   assign v3_1517448501_773 = v3_1517448501_772 & ~f125;
   assign v3_1517448501_774 = v3_1517448501_773 & ~f128;
   assign v3_1517448501_775 = v3_1517448501_774 & ~f131;
   assign v3_1517448501_776 = 1'b0; 
   assign v3_1517448501_777 = a_got_resp_initiator_2 & ~f004;
   assign v3_1517448501_779 = v3_1517448501_777 & ~f005;
   assign v3_1517448501_780 = ~v3_1517448501_781;
   assign v3_1517448501_781 = ~v3_1517448501_779 & ~f113;
   assign v3_1517448501_782 = ~v3_1517448501_783;
   assign v3_1517448501_783 = ~v3_1517448501_780 & ~f117;
   assign v3_1517448501_784 = ~v3_1517448501_785;
   assign v3_1517448501_785 = ~v3_1517448501_782 & ~f121;
   assign v3_1517448501_786 = ~v3_1517448501_787;
   assign v3_1517448501_787 = ~v3_1517448501_784 & ~f125;
   assign v3_1517448501_788 = ~v3_1517448501_789;
   assign v3_1517448501_789 = ~v3_1517448501_786 & ~f128;
   assign v3_1517448501_790 = ~v3_1517448501_791;
   assign v3_1517448501_791 = ~v3_1517448501_788 & ~f131;
   assign v3_1517448501_792 = 1'b0; 
   assign v3_1517448501_793 = ~v3_1517448501_794;
   assign v3_1517448501_794 = ~a_commited_initiator_2 & ~f004;
   assign v3_1517448501_795 = v3_1517448501_793 & ~f140;
   assign v3_1517448501_796 = v3_1517448501_795 & ~f141;
   assign v3_1517448501_797 = v3_1517448501_796 & ~f142;
   assign v3_1517448501_798 = v3_1517448501_797 & ~f143;
   assign v3_1517448501_799 = 1'b0; 
   assign v3_1517448501_800 = ~v3_1517448501_801;
   assign v3_1517448501_801 = ~a_finished_initiator_2 & ~f140;
   assign v3_1517448501_802 = ~v3_1517448501_803;
   assign v3_1517448501_803 = ~v3_1517448501_800 & ~f141;
   assign v3_1517448501_804 = ~v3_1517448501_805;
   assign v3_1517448501_805 = ~v3_1517448501_802 & ~f142;
   assign v3_1517448501_806 = ~v3_1517448501_807;
   assign v3_1517448501_807 = ~v3_1517448501_804 & ~f143;
   assign v3_1517448501_808 = 1'b0; 
   assign v3_1517448501_809 = ~v3_1517448501_810;
   assign v3_1517448501_810 = ~a_corrupted_initiator_2 & ~f005;
   assign v3_1517448501_811 = 1'b0; 
   assign v3_1517448501_812 = ~a_start_responder_0 & ~f036;
   assign v3_1517448501_813 = v3_1517448501_812 & ~f040;
   assign v3_1517448501_814 = v3_1517448501_813 & ~f044;
   assign v3_1517448501_815 = v3_1517448501_814 & ~f048;
   assign v3_1517448501_816 = v3_1517448501_815 & ~f051;
   assign v3_1517448501_817 = v3_1517448501_816 & ~f054;
   assign v3_1517448501_818 = v3_1517448501_817 & ~f057;
   assign v3_1517448501_819 = v3_1517448501_818 & ~f060;
   assign v3_1517448501_820 = v3_1517448501_819 & ~f063;
   assign v3_1517448501_821 = v3_1517448501_820 & ~f066;
   assign v3_1517448501_822 = v3_1517448501_821 & ~f069;
   assign v3_1517448501_823 = v3_1517448501_822 & ~f072;
   assign v3_1517448501_824 = v3_1517448501_823 & ~f075;
   assign v3_1517448501_825 = v3_1517448501_824 & ~f078;
   assign v3_1517448501_826 = v3_1517448501_825 & ~f081;
   assign v3_1517448501_827 = v3_1517448501_826 & ~f084;
   assign v3_1517448501_828 = v3_1517448501_827 & ~f087;
   assign v3_1517448501_829 = v3_1517448501_828 & ~f090;
   assign v3_1517448501_830 = v3_1517448501_829 & ~f093;
   assign v3_1517448501_831 = v3_1517448501_830 & ~f096;
   assign v3_1517448501_832 = v3_1517448501_831 & ~f099;
   assign v3_1517448501_833 = v3_1517448501_832 & ~f102;
   assign v3_1517448501_834 = v3_1517448501_833 & ~f105;
   assign v3_1517448501_835 = v3_1517448501_834 & ~f108;
   assign v3_1517448501_836 = 1'b0; 
   assign v3_1517448501_837 = a_got_msg_responder_0 & ~f006;
   assign v3_1517448501_839 = v3_1517448501_837 & ~f007;
   assign v3_1517448501_840 = ~v3_1517448501_841;
   assign v3_1517448501_841 = ~v3_1517448501_839 & ~f036;
   assign v3_1517448501_842 = ~v3_1517448501_843;
   assign v3_1517448501_843 = ~v3_1517448501_840 & ~f040;
   assign v3_1517448501_844 = ~v3_1517448501_845;
   assign v3_1517448501_845 = ~v3_1517448501_842 & ~f044;
   assign v3_1517448501_846 = ~v3_1517448501_847;
   assign v3_1517448501_847 = ~v3_1517448501_844 & ~f048;
   assign v3_1517448501_848 = ~v3_1517448501_849;
   assign v3_1517448501_849 = ~v3_1517448501_846 & ~f051;
   assign v3_1517448501_850 = ~v3_1517448501_851;
   assign v3_1517448501_851 = ~v3_1517448501_848 & ~f054;
   assign v3_1517448501_852 = ~v3_1517448501_853;
   assign v3_1517448501_853 = ~v3_1517448501_850 & ~f057;
   assign v3_1517448501_854 = ~v3_1517448501_855;
   assign v3_1517448501_855 = ~v3_1517448501_852 & ~f060;
   assign v3_1517448501_856 = ~v3_1517448501_857;
   assign v3_1517448501_857 = ~v3_1517448501_854 & ~f063;
   assign v3_1517448501_858 = ~v3_1517448501_859;
   assign v3_1517448501_859 = ~v3_1517448501_856 & ~f066;
   assign v3_1517448501_860 = ~v3_1517448501_861;
   assign v3_1517448501_861 = ~v3_1517448501_858 & ~f069;
   assign v3_1517448501_862 = ~v3_1517448501_863;
   assign v3_1517448501_863 = ~v3_1517448501_860 & ~f072;
   assign v3_1517448501_864 = ~v3_1517448501_865;
   assign v3_1517448501_865 = ~v3_1517448501_862 & ~f075;
   assign v3_1517448501_866 = ~v3_1517448501_867;
   assign v3_1517448501_867 = ~v3_1517448501_864 & ~f078;
   assign v3_1517448501_868 = ~v3_1517448501_869;
   assign v3_1517448501_869 = ~v3_1517448501_866 & ~f081;
   assign v3_1517448501_870 = ~v3_1517448501_871;
   assign v3_1517448501_871 = ~v3_1517448501_868 & ~f084;
   assign v3_1517448501_872 = ~v3_1517448501_873;
   assign v3_1517448501_873 = ~v3_1517448501_870 & ~f087;
   assign v3_1517448501_874 = ~v3_1517448501_875;
   assign v3_1517448501_875 = ~v3_1517448501_872 & ~f090;
   assign v3_1517448501_876 = ~v3_1517448501_877;
   assign v3_1517448501_877 = ~v3_1517448501_874 & ~f093;
   assign v3_1517448501_878 = ~v3_1517448501_879;
   assign v3_1517448501_879 = ~v3_1517448501_876 & ~f096;
   assign v3_1517448501_880 = ~v3_1517448501_881;
   assign v3_1517448501_881 = ~v3_1517448501_878 & ~f099;
   assign v3_1517448501_882 = ~v3_1517448501_883;
   assign v3_1517448501_883 = ~v3_1517448501_880 & ~f102;
   assign v3_1517448501_884 = ~v3_1517448501_885;
   assign v3_1517448501_885 = ~v3_1517448501_882 & ~f105;
   assign v3_1517448501_886 = ~v3_1517448501_887;
   assign v3_1517448501_887 = ~v3_1517448501_884 & ~f108;
   assign v3_1517448501_888 = 1'b0; 
   assign v3_1517448501_889 = ~v3_1517448501_890;
   assign v3_1517448501_890 = ~a_send_reply_responder_0 & ~f006;
   assign v3_1517448501_891 = v3_1517448501_889 & ~f111;
   assign v3_1517448501_892 = v3_1517448501_891 & ~f112;
   assign v3_1517448501_893 = v3_1517448501_892 & ~f113;
   assign v3_1517448501_894 = v3_1517448501_893 & ~f114;
   assign v3_1517448501_895 = 1'b0; 
   assign v3_1517448501_896 = ~v3_1517448501_897;
   assign v3_1517448501_897 = ~a_wait_resp_responder_0 & ~f111;
   assign v3_1517448501_898 = ~v3_1517448501_899;
   assign v3_1517448501_899 = ~v3_1517448501_896 & ~f112;
   assign v3_1517448501_900 = ~v3_1517448501_901;
   assign v3_1517448501_901 = ~v3_1517448501_898 & ~f113;
   assign v3_1517448501_902 = ~v3_1517448501_903;
   assign v3_1517448501_903 = ~v3_1517448501_900 & ~f114;
   assign v3_1517448501_904 = v3_1517448501_902 & ~f132;
   assign v3_1517448501_905 = v3_1517448501_904 & ~f136;
   assign v3_1517448501_906 = v3_1517448501_905 & ~f140;
   assign v3_1517448501_907 = v3_1517448501_906 & ~f144;
   assign v3_1517448501_908 = 1'b0; 
   assign v3_1517448501_910 = a_got_resp_responder_0 & ~f008;
   assign v3_1517448501_912 = v3_1517448501_910 & ~f009;
   assign v3_1517448501_913 = ~v3_1517448501_914;
   assign v3_1517448501_914 = ~v3_1517448501_912 & ~f132;
   assign v3_1517448501_915 = ~v3_1517448501_916;
   assign v3_1517448501_916 = ~v3_1517448501_913 & ~f136;
   assign v3_1517448501_917 = ~v3_1517448501_918;
   assign v3_1517448501_918 = ~v3_1517448501_915 & ~f140;
   assign v3_1517448501_919 = ~v3_1517448501_920;
   assign v3_1517448501_920 = ~v3_1517448501_917 & ~f144;
   assign v3_1517448501_921 = 1'b0; 
   assign v3_1517448501_922 = ~v3_1517448501_923;
   assign v3_1517448501_923 = ~a_finished_responder_0 & ~f009;
   assign v3_1517448501_924 = 1'b0; 
   assign v3_1517448501_925 = ~v3_1517448501_926;
   assign v3_1517448501_926 = ~a_corrupted_responder_0 & ~f007;
   assign v3_1517448501_927 = ~v3_1517448501_928;
   assign v3_1517448501_928 = ~v3_1517448501_925 & ~f008;
   assign v3_1517448501_929 = 1'b0; 
   assign v3_1517448501_930 = ~a_start_responder_1 & ~f037;
   assign v3_1517448501_931 = v3_1517448501_930 & ~f041;
   assign v3_1517448501_932 = v3_1517448501_931 & ~f045;
   assign v3_1517448501_933 = v3_1517448501_932 & ~f049;
   assign v3_1517448501_934 = v3_1517448501_933 & ~f052;
   assign v3_1517448501_935 = v3_1517448501_934 & ~f055;
   assign v3_1517448501_936 = v3_1517448501_935 & ~f058;
   assign v3_1517448501_937 = v3_1517448501_936 & ~f061;
   assign v3_1517448501_938 = v3_1517448501_937 & ~f064;
   assign v3_1517448501_939 = v3_1517448501_938 & ~f067;
   assign v3_1517448501_940 = v3_1517448501_939 & ~f070;
   assign v3_1517448501_941 = v3_1517448501_940 & ~f073;
   assign v3_1517448501_942 = v3_1517448501_941 & ~f076;
   assign v3_1517448501_943 = v3_1517448501_942 & ~f079;
   assign v3_1517448501_944 = v3_1517448501_943 & ~f082;
   assign v3_1517448501_945 = v3_1517448501_944 & ~f085;
   assign v3_1517448501_946 = v3_1517448501_945 & ~f088;
   assign v3_1517448501_947 = v3_1517448501_946 & ~f091;
   assign v3_1517448501_948 = v3_1517448501_947 & ~f094;
   assign v3_1517448501_949 = v3_1517448501_948 & ~f097;
   assign v3_1517448501_950 = v3_1517448501_949 & ~f100;
   assign v3_1517448501_951 = v3_1517448501_950 & ~f103;
   assign v3_1517448501_952 = v3_1517448501_951 & ~f106;
   assign v3_1517448501_953 = v3_1517448501_952 & ~f109;
   assign v3_1517448501_954 = 1'b0; 
   assign v3_1517448501_955 = a_got_msg_responder_1 & ~f010;
   assign v3_1517448501_957 = v3_1517448501_955 & ~f011;
   assign v3_1517448501_958 = ~v3_1517448501_959;
   assign v3_1517448501_959 = ~v3_1517448501_957 & ~f037;
   assign v3_1517448501_960 = ~v3_1517448501_961;
   assign v3_1517448501_961 = ~v3_1517448501_958 & ~f041;
   assign v3_1517448501_962 = ~v3_1517448501_963;
   assign v3_1517448501_963 = ~v3_1517448501_960 & ~f045;
   assign v3_1517448501_964 = ~v3_1517448501_965;
   assign v3_1517448501_965 = ~v3_1517448501_962 & ~f049;
   assign v3_1517448501_966 = ~v3_1517448501_967;
   assign v3_1517448501_967 = ~v3_1517448501_964 & ~f052;
   assign v3_1517448501_968 = ~v3_1517448501_969;
   assign v3_1517448501_969 = ~v3_1517448501_966 & ~f055;
   assign v3_1517448501_970 = ~v3_1517448501_971;
   assign v3_1517448501_971 = ~v3_1517448501_968 & ~f058;
   assign v3_1517448501_972 = ~v3_1517448501_973;
   assign v3_1517448501_973 = ~v3_1517448501_970 & ~f061;
   assign v3_1517448501_974 = ~v3_1517448501_975;
   assign v3_1517448501_975 = ~v3_1517448501_972 & ~f064;
   assign v3_1517448501_976 = ~v3_1517448501_977;
   assign v3_1517448501_977 = ~v3_1517448501_974 & ~f067;
   assign v3_1517448501_978 = ~v3_1517448501_979;
   assign v3_1517448501_979 = ~v3_1517448501_976 & ~f070;
   assign v3_1517448501_980 = ~v3_1517448501_981;
   assign v3_1517448501_981 = ~v3_1517448501_978 & ~f073;
   assign v3_1517448501_982 = ~v3_1517448501_983;
   assign v3_1517448501_983 = ~v3_1517448501_980 & ~f076;
   assign v3_1517448501_984 = ~v3_1517448501_985;
   assign v3_1517448501_985 = ~v3_1517448501_982 & ~f079;
   assign v3_1517448501_986 = ~v3_1517448501_987;
   assign v3_1517448501_987 = ~v3_1517448501_984 & ~f082;
   assign v3_1517448501_988 = ~v3_1517448501_989;
   assign v3_1517448501_989 = ~v3_1517448501_986 & ~f085;
   assign v3_1517448501_990 = ~v3_1517448501_991;
   assign v3_1517448501_991 = ~v3_1517448501_988 & ~f088;
   assign v3_1517448501_992 = ~v3_1517448501_993;
   assign v3_1517448501_993 = ~v3_1517448501_990 & ~f091;
   assign v3_1517448501_994 = ~v3_1517448501_995;
   assign v3_1517448501_995 = ~v3_1517448501_992 & ~f094;
   assign v3_1517448501_996 = ~v3_1517448501_997;
   assign v3_1517448501_997 = ~v3_1517448501_994 & ~f097;
   assign v3_1517448501_998 = ~v3_1517448501_999;
   assign v3_1517448501_999 = ~v3_1517448501_996 & ~f100;
   assign v3_1517448501_1000 = ~v3_1517448501_1001;
   assign v3_1517448501_1001 = ~v3_1517448501_998 & ~f103;
   assign v3_1517448501_1002 = ~v3_1517448501_1003;
   assign v3_1517448501_1003 = ~v3_1517448501_1000 & ~f106;
   assign v3_1517448501_1004 = ~v3_1517448501_1005;
   assign v3_1517448501_1005 = ~v3_1517448501_1002 & ~f109;
   assign v3_1517448501_1006 = 1'b0; 
   assign v3_1517448501_1007 = ~v3_1517448501_1008;
   assign v3_1517448501_1008 = ~a_send_reply_responder_1 & ~f010;
   assign v3_1517448501_1009 = v3_1517448501_1007 & ~f115;
   assign v3_1517448501_1010 = v3_1517448501_1009 & ~f116;
   assign v3_1517448501_1011 = v3_1517448501_1010 & ~f117;
   assign v3_1517448501_1012 = v3_1517448501_1011 & ~f118;
   assign v3_1517448501_1013 = 1'b0; 
   assign v3_1517448501_1014 = ~v3_1517448501_1015;
   assign v3_1517448501_1015 = ~a_wait_resp_responder_1 & ~f115;
   assign v3_1517448501_1016 = ~v3_1517448501_1017;
   assign v3_1517448501_1017 = ~v3_1517448501_1014 & ~f116;
   assign v3_1517448501_1018 = ~v3_1517448501_1019;
   assign v3_1517448501_1019 = ~v3_1517448501_1016 & ~f117;
   assign v3_1517448501_1020 = ~v3_1517448501_1021;
   assign v3_1517448501_1021 = ~v3_1517448501_1018 & ~f118;
   assign v3_1517448501_1022 = v3_1517448501_1020 & ~f133;
   assign v3_1517448501_1023 = v3_1517448501_1022 & ~f137;
   assign v3_1517448501_1024 = v3_1517448501_1023 & ~f141;
   assign v3_1517448501_1025 = v3_1517448501_1024 & ~f145;
   assign v3_1517448501_1026 = 1'b0; 
   assign v3_1517448501_1028 = a_got_resp_responder_1 & ~f012;
   assign v3_1517448501_1030 = v3_1517448501_1028 & ~f013;
   assign v3_1517448501_1031 = ~v3_1517448501_1032;
   assign v3_1517448501_1032 = ~v3_1517448501_1030 & ~f133;
   assign v3_1517448501_1033 = ~v3_1517448501_1034;
   assign v3_1517448501_1034 = ~v3_1517448501_1031 & ~f137;
   assign v3_1517448501_1035 = ~v3_1517448501_1036;
   assign v3_1517448501_1036 = ~v3_1517448501_1033 & ~f141;
   assign v3_1517448501_1037 = ~v3_1517448501_1038;
   assign v3_1517448501_1038 = ~v3_1517448501_1035 & ~f145;
   assign v3_1517448501_1039 = 1'b0; 
   assign v3_1517448501_1040 = ~v3_1517448501_1041;
   assign v3_1517448501_1041 = ~a_finished_responder_1 & ~f013;
   assign v3_1517448501_1042 = 1'b0; 
   assign v3_1517448501_1043 = ~v3_1517448501_1044;
   assign v3_1517448501_1044 = ~a_corrupted_responder_1 & ~f011;
   assign v3_1517448501_1045 = ~v3_1517448501_1046;
   assign v3_1517448501_1046 = ~v3_1517448501_1043 & ~f012;
   assign v3_1517448501_1047 = 1'b0; 
   assign v3_1517448501_1048 = ~a_start_responder_2 & ~f038;
   assign v3_1517448501_1049 = v3_1517448501_1048 & ~f042;
   assign v3_1517448501_1050 = v3_1517448501_1049 & ~f046;
   assign v3_1517448501_1051 = v3_1517448501_1050 & ~f050;
   assign v3_1517448501_1052 = v3_1517448501_1051 & ~f053;
   assign v3_1517448501_1053 = v3_1517448501_1052 & ~f056;
   assign v3_1517448501_1054 = v3_1517448501_1053 & ~f059;
   assign v3_1517448501_1055 = v3_1517448501_1054 & ~f062;
   assign v3_1517448501_1056 = v3_1517448501_1055 & ~f065;
   assign v3_1517448501_1057 = v3_1517448501_1056 & ~f068;
   assign v3_1517448501_1058 = v3_1517448501_1057 & ~f071;
   assign v3_1517448501_1059 = v3_1517448501_1058 & ~f074;
   assign v3_1517448501_1060 = v3_1517448501_1059 & ~f077;
   assign v3_1517448501_1061 = v3_1517448501_1060 & ~f080;
   assign v3_1517448501_1062 = v3_1517448501_1061 & ~f083;
   assign v3_1517448501_1063 = v3_1517448501_1062 & ~f086;
   assign v3_1517448501_1064 = v3_1517448501_1063 & ~f089;
   assign v3_1517448501_1065 = v3_1517448501_1064 & ~f092;
   assign v3_1517448501_1066 = v3_1517448501_1065 & ~f095;
   assign v3_1517448501_1067 = v3_1517448501_1066 & ~f098;
   assign v3_1517448501_1068 = v3_1517448501_1067 & ~f101;
   assign v3_1517448501_1069 = v3_1517448501_1068 & ~f104;
   assign v3_1517448501_1070 = v3_1517448501_1069 & ~f107;
   assign v3_1517448501_1071 = v3_1517448501_1070 & ~f110;
   assign v3_1517448501_1072 = 1'b0; 
   assign v3_1517448501_1073 = a_got_msg_responder_2 & ~f014;
   assign v3_1517448501_1075 = v3_1517448501_1073 & ~f015;
   assign v3_1517448501_1076 = ~v3_1517448501_1077;
   assign v3_1517448501_1077 = ~v3_1517448501_1075 & ~f038;
   assign v3_1517448501_1078 = ~v3_1517448501_1079;
   assign v3_1517448501_1079 = ~v3_1517448501_1076 & ~f042;
   assign v3_1517448501_1080 = ~v3_1517448501_1081;
   assign v3_1517448501_1081 = ~v3_1517448501_1078 & ~f046;
   assign v3_1517448501_1082 = ~v3_1517448501_1083;
   assign v3_1517448501_1083 = ~v3_1517448501_1080 & ~f050;
   assign v3_1517448501_1084 = ~v3_1517448501_1085;
   assign v3_1517448501_1085 = ~v3_1517448501_1082 & ~f053;
   assign v3_1517448501_1086 = ~v3_1517448501_1087;
   assign v3_1517448501_1087 = ~v3_1517448501_1084 & ~f056;
   assign v3_1517448501_1088 = ~v3_1517448501_1089;
   assign v3_1517448501_1089 = ~v3_1517448501_1086 & ~f059;
   assign v3_1517448501_1090 = ~v3_1517448501_1091;
   assign v3_1517448501_1091 = ~v3_1517448501_1088 & ~f062;
   assign v3_1517448501_1092 = ~v3_1517448501_1093;
   assign v3_1517448501_1093 = ~v3_1517448501_1090 & ~f065;
   assign v3_1517448501_1094 = ~v3_1517448501_1095;
   assign v3_1517448501_1095 = ~v3_1517448501_1092 & ~f068;
   assign v3_1517448501_1096 = ~v3_1517448501_1097;
   assign v3_1517448501_1097 = ~v3_1517448501_1094 & ~f071;
   assign v3_1517448501_1098 = ~v3_1517448501_1099;
   assign v3_1517448501_1099 = ~v3_1517448501_1096 & ~f074;
   assign v3_1517448501_1100 = ~v3_1517448501_1101;
   assign v3_1517448501_1101 = ~v3_1517448501_1098 & ~f077;
   assign v3_1517448501_1102 = ~v3_1517448501_1103;
   assign v3_1517448501_1103 = ~v3_1517448501_1100 & ~f080;
   assign v3_1517448501_1104 = ~v3_1517448501_1105;
   assign v3_1517448501_1105 = ~v3_1517448501_1102 & ~f083;
   assign v3_1517448501_1106 = ~v3_1517448501_1107;
   assign v3_1517448501_1107 = ~v3_1517448501_1104 & ~f086;
   assign v3_1517448501_1108 = ~v3_1517448501_1109;
   assign v3_1517448501_1109 = ~v3_1517448501_1106 & ~f089;
   assign v3_1517448501_1110 = ~v3_1517448501_1111;
   assign v3_1517448501_1111 = ~v3_1517448501_1108 & ~f092;
   assign v3_1517448501_1112 = ~v3_1517448501_1113;
   assign v3_1517448501_1113 = ~v3_1517448501_1110 & ~f095;
   assign v3_1517448501_1114 = ~v3_1517448501_1115;
   assign v3_1517448501_1115 = ~v3_1517448501_1112 & ~f098;
   assign v3_1517448501_1116 = ~v3_1517448501_1117;
   assign v3_1517448501_1117 = ~v3_1517448501_1114 & ~f101;
   assign v3_1517448501_1118 = ~v3_1517448501_1119;
   assign v3_1517448501_1119 = ~v3_1517448501_1116 & ~f104;
   assign v3_1517448501_1120 = ~v3_1517448501_1121;
   assign v3_1517448501_1121 = ~v3_1517448501_1118 & ~f107;
   assign v3_1517448501_1122 = ~v3_1517448501_1123;
   assign v3_1517448501_1123 = ~v3_1517448501_1120 & ~f110;
   assign v3_1517448501_1124 = 1'b0; 
   assign v3_1517448501_1125 = ~v3_1517448501_1126;
   assign v3_1517448501_1126 = ~a_send_reply_responder_2 & ~f014;
   assign v3_1517448501_1127 = v3_1517448501_1125 & ~f119;
   assign v3_1517448501_1128 = v3_1517448501_1127 & ~f120;
   assign v3_1517448501_1129 = v3_1517448501_1128 & ~f121;
   assign v3_1517448501_1130 = v3_1517448501_1129 & ~f122;
   assign v3_1517448501_1131 = 1'b0; 
   assign v3_1517448501_1132 = ~v3_1517448501_1133;
   assign v3_1517448501_1133 = ~a_wait_resp_responder_2 & ~f119;
   assign v3_1517448501_1134 = ~v3_1517448501_1135;
   assign v3_1517448501_1135 = ~v3_1517448501_1132 & ~f120;
   assign v3_1517448501_1136 = ~v3_1517448501_1137;
   assign v3_1517448501_1137 = ~v3_1517448501_1134 & ~f121;
   assign v3_1517448501_1138 = ~v3_1517448501_1139;
   assign v3_1517448501_1139 = ~v3_1517448501_1136 & ~f122;
   assign v3_1517448501_1140 = v3_1517448501_1138 & ~f134;
   assign v3_1517448501_1141 = v3_1517448501_1140 & ~f138;
   assign v3_1517448501_1142 = v3_1517448501_1141 & ~f142;
   assign v3_1517448501_1143 = v3_1517448501_1142 & ~f146;
   assign v3_1517448501_1144 = 1'b0; 
   assign v3_1517448501_1146 = a_got_resp_responder_2 & ~f016;
   assign v3_1517448501_1148 = v3_1517448501_1146 & ~f017;
   assign v3_1517448501_1149 = ~v3_1517448501_1150;
   assign v3_1517448501_1150 = ~v3_1517448501_1148 & ~f134;
   assign v3_1517448501_1151 = ~v3_1517448501_1152;
   assign v3_1517448501_1152 = ~v3_1517448501_1149 & ~f138;
   assign v3_1517448501_1153 = ~v3_1517448501_1154;
   assign v3_1517448501_1154 = ~v3_1517448501_1151 & ~f142;
   assign v3_1517448501_1155 = ~v3_1517448501_1156;
   assign v3_1517448501_1156 = ~v3_1517448501_1153 & ~f146;
   assign v3_1517448501_1157 = 1'b0; 
   assign v3_1517448501_1158 = ~v3_1517448501_1159;
   assign v3_1517448501_1159 = ~a_finished_responder_2 & ~f017;
   assign v3_1517448501_1160 = 1'b0; 
   assign v3_1517448501_1161 = ~v3_1517448501_1162;
   assign v3_1517448501_1162 = ~a_corrupted_responder_2 & ~f015;
   assign v3_1517448501_1163 = ~v3_1517448501_1164;
   assign v3_1517448501_1164 = ~v3_1517448501_1161 & ~f016;
   assign v3_1517448501_1165 = 1'b0; 
   assign v3_1517448501_1167 = ~v3_1517448501_1168;
   assign v3_1517448501_1168 = a_q & ~f018;
   assign v3_1517448501_1169 = ~v3_1517448501_1170;
   assign v3_1517448501_1170 = ~v3_1517448501_1167 & ~f024;
   assign v3_1517448501_1172 = ~v3_1517448501_1173;
   assign v3_1517448501_1173 = ~v3_1517448501_1169 & ~f025;
   assign v3_1517448501_1174 = ~v3_1517448501_1175;
   assign v3_1517448501_1175 = ~v3_1517448501_1172 & ~f026;
   assign v3_1517448501_1176 = ~v3_1517448501_1177;
   assign v3_1517448501_1177 = ~v3_1517448501_1174 & ~f027;
   assign v3_1517448501_1179 = ~v3_1517448501_1180;
   assign v3_1517448501_1180 = ~v3_1517448501_1176 & ~f028;
   assign v3_1517448501_1181 = ~v3_1517448501_1182;
   assign v3_1517448501_1182 = ~v3_1517448501_1179 & ~f031;
   assign v3_1517448501_1183 = ~v3_1517448501_1184;
   assign v3_1517448501_1184 = ~v3_1517448501_1181 & ~f032;
   assign v3_1517448501_1186 = ~v3_1517448501_1187;
   assign v3_1517448501_1187 = ~v3_1517448501_1183 & ~f033;
   assign v3_1517448501_1188 = ~v3_1517448501_1189;
   assign v3_1517448501_1189 = ~v3_1517448501_1186 & ~f034;
   assign v3_1517448501_1191 = ~v3_1517448501_1192;
   assign v3_1517448501_1192 = ~v3_1517448501_1188 & ~f035;
   assign v3_1517448501_1193 = v3_1517448501_1191 & ~f039;
   assign v3_1517448501_1194 = v3_1517448501_1193 & ~f043;
   assign v3_1517448501_1195 = v3_1517448501_1194 & ~f047;
   assign v3_1517448501_1196 = v3_1517448501_1195 & ~f114;
   assign v3_1517448501_1197 = v3_1517448501_1196 & ~f118;
   assign v3_1517448501_1198 = v3_1517448501_1197 & ~f122;
   assign v3_1517448501_1199 = v3_1517448501_1198 & ~f135;
   assign v3_1517448501_1200 = v3_1517448501_1199 & ~f139;
   assign v3_1517448501_1201 = v3_1517448501_1200 & ~f143;
   assign v3_1517448501_1202 = 1'b0; 
   assign v3_1517448501_1203 = a_got3 & ~f018;
   assign v3_1517448501_1205 = v3_1517448501_1203 & ~f019;
   assign v3_1517448501_1207 = v3_1517448501_1205 & ~f020;
   assign v3_1517448501_1208 = ~v3_1517448501_1209;
   assign v3_1517448501_1209 = ~v3_1517448501_1207 & ~f039;
   assign v3_1517448501_1210 = ~v3_1517448501_1211;
   assign v3_1517448501_1211 = ~v3_1517448501_1208 & ~f043;
   assign v3_1517448501_1212 = ~v3_1517448501_1213;
   assign v3_1517448501_1213 = ~v3_1517448501_1210 & ~f047;
   assign v3_1517448501_1214 = ~v3_1517448501_1215;
   assign v3_1517448501_1215 = ~v3_1517448501_1212 & ~f114;
   assign v3_1517448501_1216 = ~v3_1517448501_1217;
   assign v3_1517448501_1217 = ~v3_1517448501_1214 & ~f118;
   assign v3_1517448501_1218 = ~v3_1517448501_1219;
   assign v3_1517448501_1219 = ~v3_1517448501_1216 & ~f122;
   assign v3_1517448501_1220 = 1'b0; 
   assign v3_1517448501_1221 = ~v3_1517448501_1222;
   assign v3_1517448501_1222 = ~a_c1 & ~f019;
   assign v3_1517448501_1223 = v3_1517448501_1221 & ~f021;
   assign v3_1517448501_1224 = v3_1517448501_1223 & ~f022;
   assign v3_1517448501_1226 = v3_1517448501_1224 & ~f023;
   assign v3_1517448501_1227 = 1'b0; 
   assign v3_1517448501_1228 = ~v3_1517448501_1229;
   assign v3_1517448501_1229 = ~a_c2 & ~f021;
   assign v3_1517448501_1230 = ~v3_1517448501_1231;
   assign v3_1517448501_1231 = ~v3_1517448501_1228 & ~f022;
   assign v3_1517448501_1232 = ~v3_1517448501_1233;
   assign v3_1517448501_1233 = ~v3_1517448501_1230 & ~f023;
   assign v3_1517448501_1234 = v3_1517448501_1232 & ~f024;
   assign v3_1517448501_1235 = v3_1517448501_1234 & ~f025;
   assign v3_1517448501_1236 = 1'b0; 
   assign v3_1517448501_1237 = ~v3_1517448501_1238;
   assign v3_1517448501_1238 = ~a_d1 & ~f020;
   assign v3_1517448501_1239 = v3_1517448501_1237 & ~f026;
   assign v3_1517448501_1240 = v3_1517448501_1239 & ~f027;
   assign v3_1517448501_1241 = v3_1517448501_1240 & ~f028;
   assign v3_1517448501_1242 = 1'b0; 
   assign v3_1517448501_1244 = a_got2 & ~f029;
   assign v3_1517448501_1246 = v3_1517448501_1244 & ~f030;
   assign v3_1517448501_1247 = ~v3_1517448501_1248;
   assign v3_1517448501_1248 = ~v3_1517448501_1246 & ~f135;
   assign v3_1517448501_1249 = ~v3_1517448501_1250;
   assign v3_1517448501_1250 = ~v3_1517448501_1247 & ~f139;
   assign v3_1517448501_1251 = ~v3_1517448501_1252;
   assign v3_1517448501_1252 = ~v3_1517448501_1249 & ~f143;
   assign v3_1517448501_1253 = 1'b0; 
   assign v3_1517448501_1254 = ~v3_1517448501_1255;
   assign v3_1517448501_1255 = ~a_e1 & ~f029;
   assign v3_1517448501_1256 = v3_1517448501_1254 & ~f031;
   assign v3_1517448501_1257 = v3_1517448501_1256 & ~f032;
   assign v3_1517448501_1258 = v3_1517448501_1257 & ~f033;
   assign v3_1517448501_1259 = 1'b0; 
   assign v3_1517448501_1260 = ~v3_1517448501_1261;
   assign v3_1517448501_1261 = ~a_f1 & ~f030;
   assign v3_1517448501_1262 = v3_1517448501_1260 & ~f034;
   assign v3_1517448501_1263 = v3_1517448501_1262 & ~f035;
   assign v3_1517448501_1264 = 1'b0; 
   assign v3_1517448501_1265 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1266 = v3_1517448501_1267 ? v3_1517448501_1275 : v3_1517448501_1274;
   assign v3_1517448501_1267 = v3_1517448501_143[31];
   assign v3_1517448501_1268 = v3_1517448501_95[31];
   assign v3_1517448501_1269 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1270 = ~v3_1517448501_143 + v3_1517448501_1269;
   assign v3_1517448501_1271 = ~v3_1517448501_95 + v3_1517448501_1269;
   assign v3_1517448501_1272 = v3_1517448501_1267 ? v3_1517448501_1270 : v3_1517448501_143;
   assign v3_1517448501_1273 = v3_1517448501_1268 ? v3_1517448501_1271 : v3_1517448501_95;
   assign v3_1517448501_1274 = v3_1517448501_1272 % v3_1517448501_1273;
   assign v3_1517448501_1275 = ~v3_1517448501_1274 + v3_1517448501_1269;
   assign v3_1517448501_1276 = v3_1517448501_1265 == v3_1517448501_1266;
   assign v3_1517448501_1277 = v3_1517448501_1280 ? v3_1517448501_1287 : v3_1517448501_1286;
   assign v3_1517448501_1278 = v3_1517448501_143[31];
   assign v3_1517448501_1279 = v3_1517448501_147[31];
   assign v3_1517448501_1280 = v3_1517448501_1278 ^ v3_1517448501_1279;
   assign v3_1517448501_1281 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1282 = ~v3_1517448501_143 + v3_1517448501_1281;
   assign v3_1517448501_1283 = ~v3_1517448501_147 + v3_1517448501_1281;
   assign v3_1517448501_1284 = v3_1517448501_1278 ? v3_1517448501_1282 : v3_1517448501_143;
   assign v3_1517448501_1285 = v3_1517448501_1279 ? v3_1517448501_1283 : v3_1517448501_147;
   assign v3_1517448501_1286 = v3_1517448501_1284 / v3_1517448501_1285;
   assign v3_1517448501_1287 = ~v3_1517448501_1286 + v3_1517448501_1281;
   assign v3_1517448501_1288 = v3_1517448501_70 == v3_1517448501_1277;
   assign v3_1517448501_1289 = v3_1517448501_1276 & v3_1517448501_1288;
   assign v3_1517448501_1290 = a_got_resp_initiator_0 & v3_1517448501_1289;
   assign v3_1517448501_1291 = ~v3_1517448501_1292;
   assign v3_1517448501_1292 = f000 & ~v3_1517448501_1290;
   assign v3_1517448501_1293 = a_got_resp_initiator_0 & ~v3_1517448501_1289;
   assign v3_1517448501_1294 = ~v3_1517448501_1295;
   assign v3_1517448501_1295 = f001 & ~v3_1517448501_1293;
   assign v3_1517448501_1296 = v3_1517448501_1291 & v3_1517448501_1294;
   assign v3_1517448501_1297 = 32'b00000000_00000000_00000000_00000010; 
   assign v3_1517448501_1298 = v3_1517448501_1299 ? v3_1517448501_1307 : v3_1517448501_1306;
   assign v3_1517448501_1299 = v3_1517448501_187[31];
   assign v3_1517448501_1300 = v3_1517448501_95[31];
   assign v3_1517448501_1301 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1302 = ~v3_1517448501_187 + v3_1517448501_1301;
   assign v3_1517448501_1303 = ~v3_1517448501_95 + v3_1517448501_1301;
   assign v3_1517448501_1304 = v3_1517448501_1299 ? v3_1517448501_1302 : v3_1517448501_187;
   assign v3_1517448501_1305 = v3_1517448501_1300 ? v3_1517448501_1303 : v3_1517448501_95;
   assign v3_1517448501_1306 = v3_1517448501_1304 % v3_1517448501_1305;
   assign v3_1517448501_1307 = ~v3_1517448501_1306 + v3_1517448501_1301;
   assign v3_1517448501_1308 = v3_1517448501_1297 == v3_1517448501_1298;
   assign v3_1517448501_1309 = 32'b00000000_00000000_00000000_00001000; 
   assign v3_1517448501_1310 = v3_1517448501_1313 ? v3_1517448501_1320 : v3_1517448501_1319;
   assign v3_1517448501_1311 = v3_1517448501_187[31];
   assign v3_1517448501_1312 = v3_1517448501_147[31];
   assign v3_1517448501_1313 = v3_1517448501_1311 ^ v3_1517448501_1312;
   assign v3_1517448501_1314 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1315 = ~v3_1517448501_187 + v3_1517448501_1314;
   assign v3_1517448501_1316 = ~v3_1517448501_147 + v3_1517448501_1314;
   assign v3_1517448501_1317 = v3_1517448501_1311 ? v3_1517448501_1315 : v3_1517448501_187;
   assign v3_1517448501_1318 = v3_1517448501_1312 ? v3_1517448501_1316 : v3_1517448501_147;
   assign v3_1517448501_1319 = v3_1517448501_1317 / v3_1517448501_1318;
   assign v3_1517448501_1320 = ~v3_1517448501_1319 + v3_1517448501_1314;
   assign v3_1517448501_1321 = v3_1517448501_1309 == v3_1517448501_1310;
   assign v3_1517448501_1322 = v3_1517448501_1308 & v3_1517448501_1321;
   assign v3_1517448501_1323 = a_got_resp_initiator_1 & v3_1517448501_1322;
   assign v3_1517448501_1324 = ~v3_1517448501_1325;
   assign v3_1517448501_1325 = f002 & ~v3_1517448501_1323;
   assign v3_1517448501_1326 = v3_1517448501_1296 & v3_1517448501_1324;
   assign v3_1517448501_1327 = a_got_resp_initiator_1 & ~v3_1517448501_1322;
   assign v3_1517448501_1328 = ~v3_1517448501_1329;
   assign v3_1517448501_1329 = f003 & ~v3_1517448501_1327;
   assign v3_1517448501_1330 = v3_1517448501_1326 & v3_1517448501_1328;
   assign v3_1517448501_1331 = 32'b00000000_00000000_00000000_00000011; 
   assign v3_1517448501_1332 = v3_1517448501_1333 ? v3_1517448501_1341 : v3_1517448501_1340;
   assign v3_1517448501_1333 = v3_1517448501_230[31];
   assign v3_1517448501_1334 = v3_1517448501_95[31];
   assign v3_1517448501_1335 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1336 = ~v3_1517448501_230 + v3_1517448501_1335;
   assign v3_1517448501_1337 = ~v3_1517448501_95 + v3_1517448501_1335;
   assign v3_1517448501_1338 = v3_1517448501_1333 ? v3_1517448501_1336 : v3_1517448501_230;
   assign v3_1517448501_1339 = v3_1517448501_1334 ? v3_1517448501_1337 : v3_1517448501_95;
   assign v3_1517448501_1340 = v3_1517448501_1338 % v3_1517448501_1339;
   assign v3_1517448501_1341 = ~v3_1517448501_1340 + v3_1517448501_1335;
   assign v3_1517448501_1342 = v3_1517448501_1331 == v3_1517448501_1332;
   assign v3_1517448501_1343 = 32'b00000000_00000000_00000000_00001001; 
   assign v3_1517448501_1344 = v3_1517448501_1347 ? v3_1517448501_1354 : v3_1517448501_1353;
   assign v3_1517448501_1345 = v3_1517448501_230[31];
   assign v3_1517448501_1346 = v3_1517448501_147[31];
   assign v3_1517448501_1347 = v3_1517448501_1345 ^ v3_1517448501_1346;
   assign v3_1517448501_1348 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1349 = ~v3_1517448501_230 + v3_1517448501_1348;
   assign v3_1517448501_1350 = ~v3_1517448501_147 + v3_1517448501_1348;
   assign v3_1517448501_1351 = v3_1517448501_1345 ? v3_1517448501_1349 : v3_1517448501_230;
   assign v3_1517448501_1352 = v3_1517448501_1346 ? v3_1517448501_1350 : v3_1517448501_147;
   assign v3_1517448501_1353 = v3_1517448501_1351 / v3_1517448501_1352;
   assign v3_1517448501_1354 = ~v3_1517448501_1353 + v3_1517448501_1348;
   assign v3_1517448501_1355 = v3_1517448501_1343 == v3_1517448501_1344;
   assign v3_1517448501_1356 = v3_1517448501_1342 & v3_1517448501_1355;
   assign v3_1517448501_1357 = a_got_resp_initiator_2 & v3_1517448501_1356;
   assign v3_1517448501_1358 = ~v3_1517448501_1359;
   assign v3_1517448501_1359 = f004 & ~v3_1517448501_1357;
   assign v3_1517448501_1360 = v3_1517448501_1330 & v3_1517448501_1358;
   assign v3_1517448501_1361 = a_got_resp_initiator_2 & ~v3_1517448501_1356;
   assign v3_1517448501_1362 = ~v3_1517448501_1363;
   assign v3_1517448501_1363 = f005 & ~v3_1517448501_1361;
   assign v3_1517448501_1364 = v3_1517448501_1360 & v3_1517448501_1362;
   assign v3_1517448501_1365 = 32'b00000000_00000000_00000000_00001010; 
   assign v3_1517448501_1366 = v3_1517448501_1369 ? v3_1517448501_1376 : v3_1517448501_1375;
   assign v3_1517448501_1367 = v3_1517448501_365[31];
   assign v3_1517448501_1368 = v3_1517448501_147[31];
   assign v3_1517448501_1369 = v3_1517448501_1367 ^ v3_1517448501_1368;
   assign v3_1517448501_1370 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1371 = ~v3_1517448501_365 + v3_1517448501_1370;
   assign v3_1517448501_1372 = ~v3_1517448501_147 + v3_1517448501_1370;
   assign v3_1517448501_1373 = v3_1517448501_1367 ? v3_1517448501_1371 : v3_1517448501_365;
   assign v3_1517448501_1374 = v3_1517448501_1368 ? v3_1517448501_1372 : v3_1517448501_147;
   assign v3_1517448501_1375 = v3_1517448501_1373 / v3_1517448501_1374;
   assign v3_1517448501_1376 = ~v3_1517448501_1375 + v3_1517448501_1370;
   assign v3_1517448501_1377 = v3_1517448501_1365 == v3_1517448501_1366;
   assign v3_1517448501_1378 = a_got_msg_responder_0 & v3_1517448501_1377;
   assign v3_1517448501_1379 = ~v3_1517448501_1380;
   assign v3_1517448501_1380 = f006 & ~v3_1517448501_1378;
   assign v3_1517448501_1381 = v3_1517448501_1364 & v3_1517448501_1379;
   assign v3_1517448501_1382 = a_got_msg_responder_0 & ~v3_1517448501_1377;
   assign v3_1517448501_1383 = ~v3_1517448501_1384;
   assign v3_1517448501_1384 = f007 & ~v3_1517448501_1382;
   assign v3_1517448501_1385 = v3_1517448501_1381 & v3_1517448501_1383;
   assign v3_1517448501_1386 = 32'b00000000_00000000_00000000_00000100; 
   assign v3_1517448501_1387 = v3_1517448501_1386 == v3_1517448501_393;
   assign v3_1517448501_1388 = v3_1517448501_1365 == v3_1517448501_379;
   assign v3_1517448501_1389 = v3_1517448501_1387 & v3_1517448501_1388;
   assign v3_1517448501_1390 = a_got_resp_responder_0 & ~v3_1517448501_1389;
   assign v3_1517448501_1391 = ~v3_1517448501_1392;
   assign v3_1517448501_1392 = f008 & ~v3_1517448501_1390;
   assign v3_1517448501_1393 = v3_1517448501_1385 & v3_1517448501_1391;
   assign v3_1517448501_1394 = a_got_resp_responder_0 & v3_1517448501_1389;
   assign v3_1517448501_1395 = ~v3_1517448501_1396;
   assign v3_1517448501_1396 = f009 & ~v3_1517448501_1394;
   assign v3_1517448501_1397 = v3_1517448501_1393 & v3_1517448501_1395;
   assign v3_1517448501_1398 = 32'b00000000_00000000_00000000_00001011; 
   assign v3_1517448501_1399 = v3_1517448501_1402 ? v3_1517448501_1409 : v3_1517448501_1408;
   assign v3_1517448501_1400 = v3_1517448501_465[31];
   assign v3_1517448501_1401 = v3_1517448501_147[31];
   assign v3_1517448501_1402 = v3_1517448501_1400 ^ v3_1517448501_1401;
   assign v3_1517448501_1403 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1404 = ~v3_1517448501_465 + v3_1517448501_1403;
   assign v3_1517448501_1405 = ~v3_1517448501_147 + v3_1517448501_1403;
   assign v3_1517448501_1406 = v3_1517448501_1400 ? v3_1517448501_1404 : v3_1517448501_465;
   assign v3_1517448501_1407 = v3_1517448501_1401 ? v3_1517448501_1405 : v3_1517448501_147;
   assign v3_1517448501_1408 = v3_1517448501_1406 / v3_1517448501_1407;
   assign v3_1517448501_1409 = ~v3_1517448501_1408 + v3_1517448501_1403;
   assign v3_1517448501_1410 = v3_1517448501_1398 == v3_1517448501_1399;
   assign v3_1517448501_1411 = a_got_msg_responder_1 & v3_1517448501_1410;
   assign v3_1517448501_1412 = ~v3_1517448501_1413;
   assign v3_1517448501_1413 = f010 & ~v3_1517448501_1411;
   assign v3_1517448501_1414 = v3_1517448501_1397 & v3_1517448501_1412;
   assign v3_1517448501_1415 = a_got_msg_responder_1 & ~v3_1517448501_1410;
   assign v3_1517448501_1416 = ~v3_1517448501_1417;
   assign v3_1517448501_1417 = f011 & ~v3_1517448501_1415;
   assign v3_1517448501_1418 = v3_1517448501_1414 & v3_1517448501_1416;
   assign v3_1517448501_1419 = 32'b00000000_00000000_00000000_00000101; 
   assign v3_1517448501_1420 = v3_1517448501_1419 == v3_1517448501_493;
   assign v3_1517448501_1421 = v3_1517448501_1398 == v3_1517448501_479;
   assign v3_1517448501_1422 = v3_1517448501_1420 & v3_1517448501_1421;
   assign v3_1517448501_1423 = a_got_resp_responder_1 & ~v3_1517448501_1422;
   assign v3_1517448501_1424 = ~v3_1517448501_1425;
   assign v3_1517448501_1425 = f012 & ~v3_1517448501_1423;
   assign v3_1517448501_1426 = v3_1517448501_1418 & v3_1517448501_1424;
   assign v3_1517448501_1427 = a_got_resp_responder_1 & v3_1517448501_1422;
   assign v3_1517448501_1428 = ~v3_1517448501_1429;
   assign v3_1517448501_1429 = f013 & ~v3_1517448501_1427;
   assign v3_1517448501_1430 = v3_1517448501_1426 & v3_1517448501_1428;
   assign v3_1517448501_1431 = 32'b00000000_00000000_00000000_00001100; 
   assign v3_1517448501_1432 = v3_1517448501_1435 ? v3_1517448501_1442 : v3_1517448501_1441;
   assign v3_1517448501_1433 = v3_1517448501_565[31];
   assign v3_1517448501_1434 = v3_1517448501_147[31];
   assign v3_1517448501_1435 = v3_1517448501_1433 ^ v3_1517448501_1434;
   assign v3_1517448501_1436 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1437 = ~v3_1517448501_565 + v3_1517448501_1436;
   assign v3_1517448501_1438 = ~v3_1517448501_147 + v3_1517448501_1436;
   assign v3_1517448501_1439 = v3_1517448501_1433 ? v3_1517448501_1437 : v3_1517448501_565;
   assign v3_1517448501_1440 = v3_1517448501_1434 ? v3_1517448501_1438 : v3_1517448501_147;
   assign v3_1517448501_1441 = v3_1517448501_1439 / v3_1517448501_1440;
   assign v3_1517448501_1442 = ~v3_1517448501_1441 + v3_1517448501_1436;
   assign v3_1517448501_1443 = v3_1517448501_1431 == v3_1517448501_1432;
   assign v3_1517448501_1444 = a_got_msg_responder_2 & v3_1517448501_1443;
   assign v3_1517448501_1445 = ~v3_1517448501_1446;
   assign v3_1517448501_1446 = f014 & ~v3_1517448501_1444;
   assign v3_1517448501_1447 = v3_1517448501_1430 & v3_1517448501_1445;
   assign v3_1517448501_1448 = a_got_msg_responder_2 & ~v3_1517448501_1443;
   assign v3_1517448501_1449 = ~v3_1517448501_1450;
   assign v3_1517448501_1450 = f015 & ~v3_1517448501_1448;
   assign v3_1517448501_1451 = v3_1517448501_1447 & v3_1517448501_1449;
   assign v3_1517448501_1452 = 32'b00000000_00000000_00000000_00000110; 
   assign v3_1517448501_1453 = v3_1517448501_1452 == v3_1517448501_593;
   assign v3_1517448501_1454 = v3_1517448501_1431 == v3_1517448501_579;
   assign v3_1517448501_1455 = v3_1517448501_1453 & v3_1517448501_1454;
   assign v3_1517448501_1456 = a_got_resp_responder_2 & ~v3_1517448501_1455;
   assign v3_1517448501_1457 = ~v3_1517448501_1458;
   assign v3_1517448501_1458 = f016 & ~v3_1517448501_1456;
   assign v3_1517448501_1459 = v3_1517448501_1451 & v3_1517448501_1457;
   assign v3_1517448501_1460 = a_got_resp_responder_2 & v3_1517448501_1455;
   assign v3_1517448501_1461 = ~v3_1517448501_1462;
   assign v3_1517448501_1462 = f017 & ~v3_1517448501_1460;
   assign v3_1517448501_1463 = v3_1517448501_1459 & v3_1517448501_1461;
   assign v3_1517448501_1464 = ~v3_1517448501_1465;
   assign v3_1517448501_1465 = ~a_got3 & f018;
   assign v3_1517448501_1466 = v3_1517448501_1463 & v3_1517448501_1464;
   assign v3_1517448501_1467 = {v_m_intruder, v3_1517448501_71};
   assign v3_1517448501_1468 = v3_1517448501_1471 ? ~v3_1517448501_1470 : v3_1517448501_1469;
   assign v3_1517448501_1469 = v3_1517448501_1467 >> v3_1517448501_73;
   assign v3_1517448501_1470 = ~v3_1517448501_1467 >> v3_1517448501_73;
   assign v3_1517448501_1471 = v3_1517448501_1467[31];
   assign v3_1517448501_1472 = v3_1517448501_1475 ? v3_1517448501_1482 : v3_1517448501_1481;
   assign v3_1517448501_1473 = v3_1517448501_1468[31];
   assign v3_1517448501_1474 = v3_1517448501_147[31];
   assign v3_1517448501_1475 = v3_1517448501_1473 ^ v3_1517448501_1474;
   assign v3_1517448501_1476 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1477 = ~v3_1517448501_1468 + v3_1517448501_1476;
   assign v3_1517448501_1478 = ~v3_1517448501_147 + v3_1517448501_1476;
   assign v3_1517448501_1479 = v3_1517448501_1473 ? v3_1517448501_1477 : v3_1517448501_1468;
   assign v3_1517448501_1480 = v3_1517448501_1474 ? v3_1517448501_1478 : v3_1517448501_147;
   assign v3_1517448501_1481 = v3_1517448501_1479 / v3_1517448501_1480;
   assign v3_1517448501_1482 = ~v3_1517448501_1481 + v3_1517448501_1476;
   assign v3_1517448501_1483 = v3_1517448501_1331 == v3_1517448501_1472;
   assign v3_1517448501_1484 = a_got3 & v3_1517448501_1483;
   assign v3_1517448501_1485 = ~v3_1517448501_1486;
   assign v3_1517448501_1486 = f019 & ~v3_1517448501_1484;
   assign v3_1517448501_1487 = v3_1517448501_1466 & v3_1517448501_1485;
   assign v3_1517448501_1488 = a_got3 & ~v3_1517448501_1483;
   assign v3_1517448501_1489 = ~v3_1517448501_1490;
   assign v3_1517448501_1490 = f020 & ~v3_1517448501_1488;
   assign v3_1517448501_1491 = v3_1517448501_1487 & v3_1517448501_1489;
   assign v3_1517448501_1492 = v3_1517448501_1493 ? v3_1517448501_1501 : v3_1517448501_1500;
   assign v3_1517448501_1493 = v3_1517448501_1468[31];
   assign v3_1517448501_1494 = v3_1517448501_95[31];
   assign v3_1517448501_1495 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1496 = ~v3_1517448501_1468 + v3_1517448501_1495;
   assign v3_1517448501_1497 = ~v3_1517448501_95 + v3_1517448501_1495;
   assign v3_1517448501_1498 = v3_1517448501_1493 ? v3_1517448501_1496 : v3_1517448501_1468;
   assign v3_1517448501_1499 = v3_1517448501_1494 ? v3_1517448501_1497 : v3_1517448501_95;
   assign v3_1517448501_1500 = v3_1517448501_1498 % v3_1517448501_1499;
   assign v3_1517448501_1501 = ~v3_1517448501_1500 + v3_1517448501_1495;
   assign v3_1517448501_1502 = v3_1517448501_1265 == v3_1517448501_1492;
   assign v3_1517448501_1503 = a_c1 & v3_1517448501_1502;
   assign v3_1517448501_1504 = ~v3_1517448501_1505;
   assign v3_1517448501_1505 = f021 & ~v3_1517448501_1503;
   assign v3_1517448501_1506 = v3_1517448501_1491 & v3_1517448501_1504;
   assign v3_1517448501_1507 = v3_1517448501_1386 == v3_1517448501_1492;
   assign v3_1517448501_1508 = a_c1 & v3_1517448501_1507;
   assign v3_1517448501_1509 = ~v3_1517448501_1510;
   assign v3_1517448501_1510 = f022 & ~v3_1517448501_1508;
   assign v3_1517448501_1511 = v3_1517448501_1506 & v3_1517448501_1509;
   assign v3_1517448501_1512 = ~v3_1517448501_1502 & ~v3_1517448501_1507;
   assign v3_1517448501_1513 = a_c1 & v3_1517448501_1512;
   assign v3_1517448501_1514 = ~v3_1517448501_1515;
   assign v3_1517448501_1515 = f023 & ~v3_1517448501_1513;
   assign v3_1517448501_1516 = v3_1517448501_1511 & v3_1517448501_1514;
   assign v3_1517448501_1517 = v3_1517448501_1518 ? v3_1517448501_1526 : v3_1517448501_1525;
   assign v3_1517448501_1518 = v3_1517448501_1468[31];
   assign v3_1517448501_1519 = v3_1517448501_147[31];
   assign v3_1517448501_1520 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1521 = ~v3_1517448501_1468 + v3_1517448501_1520;
   assign v3_1517448501_1522 = ~v3_1517448501_147 + v3_1517448501_1520;
   assign v3_1517448501_1523 = v3_1517448501_1518 ? v3_1517448501_1521 : v3_1517448501_1468;
   assign v3_1517448501_1524 = v3_1517448501_1519 ? v3_1517448501_1522 : v3_1517448501_147;
   assign v3_1517448501_1525 = v3_1517448501_1523 % v3_1517448501_1524;
   assign v3_1517448501_1526 = ~v3_1517448501_1525 + v3_1517448501_1520;
   assign v3_1517448501_1527 = v3_1517448501_1530 ? v3_1517448501_1537 : v3_1517448501_1536;
   assign v3_1517448501_1528 = v3_1517448501_1517[31];
   assign v3_1517448501_1529 = v3_1517448501_95[31];
   assign v3_1517448501_1530 = v3_1517448501_1528 ^ v3_1517448501_1529;
   assign v3_1517448501_1531 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1532 = ~v3_1517448501_1517 + v3_1517448501_1531;
   assign v3_1517448501_1533 = ~v3_1517448501_95 + v3_1517448501_1531;
   assign v3_1517448501_1534 = v3_1517448501_1528 ? v3_1517448501_1532 : v3_1517448501_1517;
   assign v3_1517448501_1535 = v3_1517448501_1529 ? v3_1517448501_1533 : v3_1517448501_95;
   assign v3_1517448501_1536 = v3_1517448501_1534 / v3_1517448501_1535;
   assign v3_1517448501_1537 = ~v3_1517448501_1536 + v3_1517448501_1531;
   assign v3_1517448501_1538 = v3_1517448501_1365 == v3_1517448501_1527;
   assign v3_1517448501_1539 = v3_1517448501_1507 & v3_1517448501_1538;
   assign v3_1517448501_1540 = a_c2 & v3_1517448501_1539;
   assign v3_1517448501_1541 = ~v3_1517448501_1542;
   assign v3_1517448501_1542 = f024 & ~v3_1517448501_1540;
   assign v3_1517448501_1543 = v3_1517448501_1516 & v3_1517448501_1541;
   assign v3_1517448501_1544 = a_c2 & ~v3_1517448501_1539;
   assign v3_1517448501_1545 = ~v3_1517448501_1546;
   assign v3_1517448501_1546 = f025 & ~v3_1517448501_1544;
   assign v3_1517448501_1547 = v3_1517448501_1543 & v3_1517448501_1545;
   assign v3_1517448501_1548 = v3_1517448501_70 == v3_1517448501_1527;
   assign v3_1517448501_1549 = v3_1517448501_1502 & v3_1517448501_1548;
   assign v3_1517448501_1550 = v3_1517448501_1365 == v3_1517448501_1472;
   assign v3_1517448501_1551 = v3_1517448501_1549 & v3_1517448501_1550;
   assign v3_1517448501_1552 = a_d1 & v3_1517448501_1551;
   assign v3_1517448501_1553 = ~v3_1517448501_1554;
   assign v3_1517448501_1554 = f026 & ~v3_1517448501_1552;
   assign v3_1517448501_1555 = v3_1517448501_1547 & v3_1517448501_1553;
   assign v3_1517448501_1556 = v3_1517448501_1386 == v3_1517448501_1527;
   assign v3_1517448501_1557 = v3_1517448501_1502 & v3_1517448501_1556;
   assign v3_1517448501_1558 = v3_1517448501_70 == v3_1517448501_1472;
   assign v3_1517448501_1559 = v3_1517448501_1557 & v3_1517448501_1558;
   assign v3_1517448501_1560 = a_d1 & v3_1517448501_1559;
   assign v3_1517448501_1561 = ~v3_1517448501_1562;
   assign v3_1517448501_1562 = f027 & ~v3_1517448501_1560;
   assign v3_1517448501_1563 = v3_1517448501_1555 & v3_1517448501_1561;
   assign v3_1517448501_1564 = ~v3_1517448501_1565;
   assign v3_1517448501_1565 = ~a_d1 & f028;
   assign v3_1517448501_1566 = v3_1517448501_1563 & v3_1517448501_1564;
   assign v3_1517448501_1567 = v3_1517448501_1331 == v3_1517448501_1527;
   assign v3_1517448501_1568 = a_got2 & v3_1517448501_1567;
   assign v3_1517448501_1569 = ~v3_1517448501_1570;
   assign v3_1517448501_1570 = f029 & ~v3_1517448501_1568;
   assign v3_1517448501_1571 = v3_1517448501_1566 & v3_1517448501_1569;
   assign v3_1517448501_1572 = a_got2 & ~v3_1517448501_1567;
   assign v3_1517448501_1573 = ~v3_1517448501_1574;
   assign v3_1517448501_1574 = f030 & ~v3_1517448501_1572;
   assign v3_1517448501_1575 = v3_1517448501_1571 & v3_1517448501_1573;
   assign v3_1517448501_1576 = a_e1 & v3_1517448501_1502;
   assign v3_1517448501_1577 = ~v3_1517448501_1578;
   assign v3_1517448501_1578 = f031 & ~v3_1517448501_1576;
   assign v3_1517448501_1579 = v3_1517448501_1575 & v3_1517448501_1577;
   assign v3_1517448501_1580 = a_e1 & v3_1517448501_1507;
   assign v3_1517448501_1581 = ~v3_1517448501_1582;
   assign v3_1517448501_1582 = f032 & ~v3_1517448501_1580;
   assign v3_1517448501_1583 = v3_1517448501_1579 & v3_1517448501_1581;
   assign v3_1517448501_1584 = a_e1 & v3_1517448501_1512;
   assign v3_1517448501_1585 = ~v3_1517448501_1586;
   assign v3_1517448501_1586 = f033 & ~v3_1517448501_1584;
   assign v3_1517448501_1587 = v3_1517448501_1583 & v3_1517448501_1585;
   assign v3_1517448501_1588 = a_f1 & v3_1517448501_1539;
   assign v3_1517448501_1589 = ~v3_1517448501_1590;
   assign v3_1517448501_1590 = f034 & ~v3_1517448501_1588;
   assign v3_1517448501_1591 = v3_1517448501_1587 & v3_1517448501_1589;
   assign v3_1517448501_1592 = a_f1 & ~v3_1517448501_1539;
   assign v3_1517448501_1593 = ~v3_1517448501_1594;
   assign v3_1517448501_1594 = f035 & ~v3_1517448501_1592;
   assign v3_1517448501_1595 = v3_1517448501_1591 & v3_1517448501_1593;
   assign v3_1517448501_1596 = ~a_start_initiator_0 & ~a_start_responder_0;
   assign v3_1517448501_1597 = ~v3_1517448501_1598;
   assign v3_1517448501_1598 = f036 & ~v3_1517448501_1596;
   assign v3_1517448501_1599 = v3_1517448501_1595 & v3_1517448501_1597;
   assign v3_1517448501_1600 = ~a_start_initiator_0 & ~a_start_responder_1;
   assign v3_1517448501_1601 = ~v3_1517448501_1602;
   assign v3_1517448501_1602 = f037 & ~v3_1517448501_1600;
   assign v3_1517448501_1603 = v3_1517448501_1599 & v3_1517448501_1601;
   assign v3_1517448501_1604 = ~a_start_initiator_0 & ~a_start_responder_2;
   assign v3_1517448501_1605 = ~v3_1517448501_1606;
   assign v3_1517448501_1606 = f038 & ~v3_1517448501_1604;
   assign v3_1517448501_1607 = v3_1517448501_1603 & v3_1517448501_1605;
   assign v3_1517448501_1608 = ~a_start_initiator_0 & ~a_q;
   assign v3_1517448501_1609 = ~v3_1517448501_1610;
   assign v3_1517448501_1610 = f039 & ~v3_1517448501_1608;
   assign v3_1517448501_1611 = v3_1517448501_1607 & v3_1517448501_1609;
   assign v3_1517448501_1612 = ~a_start_initiator_1 & ~a_start_responder_0;
   assign v3_1517448501_1613 = ~v3_1517448501_1614;
   assign v3_1517448501_1614 = f040 & ~v3_1517448501_1612;
   assign v3_1517448501_1615 = v3_1517448501_1611 & v3_1517448501_1613;
   assign v3_1517448501_1616 = ~a_start_initiator_1 & ~a_start_responder_1;
   assign v3_1517448501_1617 = ~v3_1517448501_1618;
   assign v3_1517448501_1618 = f041 & ~v3_1517448501_1616;
   assign v3_1517448501_1619 = v3_1517448501_1615 & v3_1517448501_1617;
   assign v3_1517448501_1620 = ~a_start_initiator_1 & ~a_start_responder_2;
   assign v3_1517448501_1621 = ~v3_1517448501_1622;
   assign v3_1517448501_1622 = f042 & ~v3_1517448501_1620;
   assign v3_1517448501_1623 = v3_1517448501_1619 & v3_1517448501_1621;
   assign v3_1517448501_1624 = ~a_start_initiator_1 & ~a_q;
   assign v3_1517448501_1625 = ~v3_1517448501_1626;
   assign v3_1517448501_1626 = f043 & ~v3_1517448501_1624;
   assign v3_1517448501_1627 = v3_1517448501_1623 & v3_1517448501_1625;
   assign v3_1517448501_1628 = ~a_start_initiator_2 & ~a_start_responder_0;
   assign v3_1517448501_1629 = ~v3_1517448501_1630;
   assign v3_1517448501_1630 = f044 & ~v3_1517448501_1628;
   assign v3_1517448501_1631 = v3_1517448501_1627 & v3_1517448501_1629;
   assign v3_1517448501_1632 = ~a_start_initiator_2 & ~a_start_responder_1;
   assign v3_1517448501_1633 = ~v3_1517448501_1634;
   assign v3_1517448501_1634 = f045 & ~v3_1517448501_1632;
   assign v3_1517448501_1635 = v3_1517448501_1631 & v3_1517448501_1633;
   assign v3_1517448501_1636 = ~a_start_initiator_2 & ~a_start_responder_2;
   assign v3_1517448501_1637 = ~v3_1517448501_1638;
   assign v3_1517448501_1638 = f046 & ~v3_1517448501_1636;
   assign v3_1517448501_1639 = v3_1517448501_1635 & v3_1517448501_1637;
   assign v3_1517448501_1640 = ~a_start_initiator_2 & ~a_q;
   assign v3_1517448501_1641 = ~v3_1517448501_1642;
   assign v3_1517448501_1642 = f047 & ~v3_1517448501_1640;
   assign v3_1517448501_1643 = v3_1517448501_1639 & v3_1517448501_1641;
   assign v3_1517448501_1644 = ~a_start_responder_0 & ~a_q;
   assign v3_1517448501_1645 = ~v3_1517448501_1646;
   assign v3_1517448501_1646 = f048 & ~v3_1517448501_1644;
   assign v3_1517448501_1647 = v3_1517448501_1643 & v3_1517448501_1645;
   assign v3_1517448501_1648 = ~a_start_responder_1 & ~a_q;
   assign v3_1517448501_1649 = ~v3_1517448501_1650;
   assign v3_1517448501_1650 = f049 & ~v3_1517448501_1648;
   assign v3_1517448501_1651 = v3_1517448501_1647 & v3_1517448501_1649;
   assign v3_1517448501_1652 = ~a_start_responder_2 & ~a_q;
   assign v3_1517448501_1653 = ~v3_1517448501_1654;
   assign v3_1517448501_1654 = f050 & ~v3_1517448501_1652;
   assign v3_1517448501_1655 = v3_1517448501_1651 & v3_1517448501_1653;
   assign v3_1517448501_1656 = ~v3_1517448501_1657;
   assign v3_1517448501_1657 = ~v3_1517448501_1644 & f051;
   assign v3_1517448501_1658 = v3_1517448501_1655 & v3_1517448501_1656;
   assign v3_1517448501_1659 = ~v3_1517448501_1660;
   assign v3_1517448501_1660 = ~v3_1517448501_1648 & f052;
   assign v3_1517448501_1661 = v3_1517448501_1658 & v3_1517448501_1659;
   assign v3_1517448501_1662 = ~v3_1517448501_1663;
   assign v3_1517448501_1663 = ~v3_1517448501_1652 & f053;
   assign v3_1517448501_1664 = v3_1517448501_1661 & v3_1517448501_1662;
   assign v3_1517448501_1665 = ~v3_1517448501_1666;
   assign v3_1517448501_1666 = ~v3_1517448501_1644 & f054;
   assign v3_1517448501_1667 = v3_1517448501_1664 & v3_1517448501_1665;
   assign v3_1517448501_1668 = ~v3_1517448501_1669;
   assign v3_1517448501_1669 = ~v3_1517448501_1648 & f055;
   assign v3_1517448501_1670 = v3_1517448501_1667 & v3_1517448501_1668;
   assign v3_1517448501_1671 = ~v3_1517448501_1672;
   assign v3_1517448501_1672 = ~v3_1517448501_1652 & f056;
   assign v3_1517448501_1673 = v3_1517448501_1670 & v3_1517448501_1671;
   assign v3_1517448501_1674 = ~v3_1517448501_1675;
   assign v3_1517448501_1675 = ~v3_1517448501_1644 & f057;
   assign v3_1517448501_1676 = v3_1517448501_1673 & v3_1517448501_1674;
   assign v3_1517448501_1677 = ~v3_1517448501_1678;
   assign v3_1517448501_1678 = ~v3_1517448501_1648 & f058;
   assign v3_1517448501_1679 = v3_1517448501_1676 & v3_1517448501_1677;
   assign v3_1517448501_1680 = ~v3_1517448501_1681;
   assign v3_1517448501_1681 = ~v3_1517448501_1652 & f059;
   assign v3_1517448501_1682 = v3_1517448501_1679 & v3_1517448501_1680;
   assign v3_1517448501_1683 = ~v3_1517448501_1684;
   assign v3_1517448501_1684 = ~v3_1517448501_1644 & f060;
   assign v3_1517448501_1685 = v3_1517448501_1682 & v3_1517448501_1683;
   assign v3_1517448501_1686 = ~v3_1517448501_1687;
   assign v3_1517448501_1687 = ~v3_1517448501_1648 & f061;
   assign v3_1517448501_1688 = v3_1517448501_1685 & v3_1517448501_1686;
   assign v3_1517448501_1689 = ~v3_1517448501_1690;
   assign v3_1517448501_1690 = ~v3_1517448501_1652 & f062;
   assign v3_1517448501_1691 = v3_1517448501_1688 & v3_1517448501_1689;
   assign v3_1517448501_1692 = ~v3_1517448501_1693;
   assign v3_1517448501_1693 = ~v3_1517448501_1644 & f063;
   assign v3_1517448501_1694 = v3_1517448501_1691 & v3_1517448501_1692;
   assign v3_1517448501_1695 = ~v3_1517448501_1696;
   assign v3_1517448501_1696 = ~v3_1517448501_1648 & f064;
   assign v3_1517448501_1697 = v3_1517448501_1694 & v3_1517448501_1695;
   assign v3_1517448501_1698 = ~v3_1517448501_1699;
   assign v3_1517448501_1699 = ~v3_1517448501_1652 & f065;
   assign v3_1517448501_1700 = v3_1517448501_1697 & v3_1517448501_1698;
   assign v3_1517448501_1701 = ~v3_1517448501_1702;
   assign v3_1517448501_1702 = ~v3_1517448501_1644 & f066;
   assign v3_1517448501_1703 = v3_1517448501_1700 & v3_1517448501_1701;
   assign v3_1517448501_1704 = ~v3_1517448501_1705;
   assign v3_1517448501_1705 = ~v3_1517448501_1648 & f067;
   assign v3_1517448501_1706 = v3_1517448501_1703 & v3_1517448501_1704;
   assign v3_1517448501_1707 = ~v3_1517448501_1708;
   assign v3_1517448501_1708 = ~v3_1517448501_1652 & f068;
   assign v3_1517448501_1709 = v3_1517448501_1706 & v3_1517448501_1707;
   assign v3_1517448501_1710 = ~v3_1517448501_1711;
   assign v3_1517448501_1711 = ~v3_1517448501_1644 & f069;
   assign v3_1517448501_1712 = v3_1517448501_1709 & v3_1517448501_1710;
   assign v3_1517448501_1713 = ~v3_1517448501_1714;
   assign v3_1517448501_1714 = ~v3_1517448501_1648 & f070;
   assign v3_1517448501_1715 = v3_1517448501_1712 & v3_1517448501_1713;
   assign v3_1517448501_1716 = ~v3_1517448501_1717;
   assign v3_1517448501_1717 = ~v3_1517448501_1652 & f071;
   assign v3_1517448501_1718 = v3_1517448501_1715 & v3_1517448501_1716;
   assign v3_1517448501_1719 = ~v3_1517448501_1720;
   assign v3_1517448501_1720 = ~v3_1517448501_1644 & f072;
   assign v3_1517448501_1721 = v3_1517448501_1718 & v3_1517448501_1719;
   assign v3_1517448501_1722 = ~v3_1517448501_1723;
   assign v3_1517448501_1723 = ~v3_1517448501_1648 & f073;
   assign v3_1517448501_1724 = v3_1517448501_1721 & v3_1517448501_1722;
   assign v3_1517448501_1725 = ~v3_1517448501_1726;
   assign v3_1517448501_1726 = ~v3_1517448501_1652 & f074;
   assign v3_1517448501_1727 = v3_1517448501_1724 & v3_1517448501_1725;
   assign v3_1517448501_1728 = ~v3_1517448501_1729;
   assign v3_1517448501_1729 = ~v3_1517448501_1644 & f075;
   assign v3_1517448501_1730 = v3_1517448501_1727 & v3_1517448501_1728;
   assign v3_1517448501_1731 = ~v3_1517448501_1732;
   assign v3_1517448501_1732 = ~v3_1517448501_1648 & f076;
   assign v3_1517448501_1733 = v3_1517448501_1730 & v3_1517448501_1731;
   assign v3_1517448501_1734 = ~v3_1517448501_1735;
   assign v3_1517448501_1735 = ~v3_1517448501_1652 & f077;
   assign v3_1517448501_1736 = v3_1517448501_1733 & v3_1517448501_1734;
   assign v3_1517448501_1737 = ~v3_1517448501_1738;
   assign v3_1517448501_1738 = ~v3_1517448501_1644 & f078;
   assign v3_1517448501_1739 = v3_1517448501_1736 & v3_1517448501_1737;
   assign v3_1517448501_1740 = ~v3_1517448501_1741;
   assign v3_1517448501_1741 = ~v3_1517448501_1648 & f079;
   assign v3_1517448501_1742 = v3_1517448501_1739 & v3_1517448501_1740;
   assign v3_1517448501_1743 = ~v3_1517448501_1744;
   assign v3_1517448501_1744 = ~v3_1517448501_1652 & f080;
   assign v3_1517448501_1745 = v3_1517448501_1742 & v3_1517448501_1743;
   assign v3_1517448501_1746 = ~v3_1517448501_1747;
   assign v3_1517448501_1747 = ~v3_1517448501_1644 & f081;
   assign v3_1517448501_1748 = v3_1517448501_1745 & v3_1517448501_1746;
   assign v3_1517448501_1749 = ~v3_1517448501_1750;
   assign v3_1517448501_1750 = ~v3_1517448501_1648 & f082;
   assign v3_1517448501_1751 = v3_1517448501_1748 & v3_1517448501_1749;
   assign v3_1517448501_1752 = ~v3_1517448501_1753;
   assign v3_1517448501_1753 = ~v3_1517448501_1652 & f083;
   assign v3_1517448501_1754 = v3_1517448501_1751 & v3_1517448501_1752;
   assign v3_1517448501_1755 = ~a_start_responder_0 & ~a_q;
   assign v3_1517448501_1756 = v3_1517448501_607 == v_kNa;
   assign v3_1517448501_1757 = v3_1517448501_1755 & v3_1517448501_1756;
   assign v3_1517448501_1758 = ~v3_1517448501_1759;
   assign v3_1517448501_1759 = f084 & ~v3_1517448501_1757;
   assign v3_1517448501_1760 = v3_1517448501_1754 & v3_1517448501_1758;
   assign v3_1517448501_1761 = ~a_start_responder_1 & ~a_q;
   assign v3_1517448501_1762 = v3_1517448501_1761 & v3_1517448501_1756;
   assign v3_1517448501_1763 = ~v3_1517448501_1764;
   assign v3_1517448501_1764 = f085 & ~v3_1517448501_1762;
   assign v3_1517448501_1765 = v3_1517448501_1760 & v3_1517448501_1763;
   assign v3_1517448501_1766 = ~a_start_responder_2 & ~a_q;
   assign v3_1517448501_1767 = v3_1517448501_1766 & v3_1517448501_1756;
   assign v3_1517448501_1768 = ~v3_1517448501_1769;
   assign v3_1517448501_1769 = f086 & ~v3_1517448501_1767;
   assign v3_1517448501_1770 = v3_1517448501_1765 & v3_1517448501_1768;
   assign v3_1517448501_1771 = ~v3_1517448501_1772;
   assign v3_1517448501_1772 = ~v3_1517448501_1757 & f087;
   assign v3_1517448501_1773 = v3_1517448501_1770 & v3_1517448501_1771;
   assign v3_1517448501_1774 = ~v3_1517448501_1775;
   assign v3_1517448501_1775 = ~v3_1517448501_1762 & f088;
   assign v3_1517448501_1776 = v3_1517448501_1773 & v3_1517448501_1774;
   assign v3_1517448501_1777 = ~v3_1517448501_1778;
   assign v3_1517448501_1778 = ~v3_1517448501_1767 & f089;
   assign v3_1517448501_1779 = v3_1517448501_1776 & v3_1517448501_1777;
   assign v3_1517448501_1780 = ~v3_1517448501_1781;
   assign v3_1517448501_1781 = ~v3_1517448501_1757 & f090;
   assign v3_1517448501_1782 = v3_1517448501_1779 & v3_1517448501_1780;
   assign v3_1517448501_1783 = ~v3_1517448501_1784;
   assign v3_1517448501_1784 = ~v3_1517448501_1762 & f091;
   assign v3_1517448501_1785 = v3_1517448501_1782 & v3_1517448501_1783;
   assign v3_1517448501_1786 = ~v3_1517448501_1787;
   assign v3_1517448501_1787 = ~v3_1517448501_1767 & f092;
   assign v3_1517448501_1788 = v3_1517448501_1785 & v3_1517448501_1786;
   assign v3_1517448501_1789 = ~a_start_responder_0 & ~a_q;
   assign v3_1517448501_1790 = 8'b00000000; 
   assign v3_1517448501_1791 = v3_1517448501_1790 == v_k_Na_A__B;
   assign v3_1517448501_1792 = ~v3_1517448501_1793;
   assign v3_1517448501_1793 = ~v3_1517448501_1756 & v3_1517448501_1791;
   assign v3_1517448501_1794 = v3_1517448501_1789 & v3_1517448501_1792;
   assign v3_1517448501_1795 = ~v3_1517448501_1796;
   assign v3_1517448501_1796 = f093 & ~v3_1517448501_1794;
   assign v3_1517448501_1797 = v3_1517448501_1788 & v3_1517448501_1795;
   assign v3_1517448501_1798 = ~a_start_responder_1 & ~a_q;
   assign v3_1517448501_1799 = v3_1517448501_1798 & v3_1517448501_1792;
   assign v3_1517448501_1800 = ~v3_1517448501_1801;
   assign v3_1517448501_1801 = f094 & ~v3_1517448501_1799;
   assign v3_1517448501_1802 = v3_1517448501_1797 & v3_1517448501_1800;
   assign v3_1517448501_1803 = ~a_start_responder_2 & ~a_q;
   assign v3_1517448501_1804 = v3_1517448501_1803 & v3_1517448501_1792;
   assign v3_1517448501_1805 = ~v3_1517448501_1806;
   assign v3_1517448501_1806 = f095 & ~v3_1517448501_1804;
   assign v3_1517448501_1807 = v3_1517448501_1802 & v3_1517448501_1805;
   assign v3_1517448501_1808 = ~v3_1517448501_1809;
   assign v3_1517448501_1809 = ~v3_1517448501_1757 & f096;
   assign v3_1517448501_1810 = v3_1517448501_1807 & v3_1517448501_1808;
   assign v3_1517448501_1811 = ~v3_1517448501_1812;
   assign v3_1517448501_1812 = ~v3_1517448501_1762 & f097;
   assign v3_1517448501_1813 = v3_1517448501_1810 & v3_1517448501_1811;
   assign v3_1517448501_1814 = ~v3_1517448501_1815;
   assign v3_1517448501_1815 = ~v3_1517448501_1767 & f098;
   assign v3_1517448501_1816 = v3_1517448501_1813 & v3_1517448501_1814;
   assign v3_1517448501_1817 = ~v3_1517448501_1818;
   assign v3_1517448501_1818 = ~v3_1517448501_1757 & f099;
   assign v3_1517448501_1819 = v3_1517448501_1816 & v3_1517448501_1817;
   assign v3_1517448501_1820 = ~v3_1517448501_1821;
   assign v3_1517448501_1821 = ~v3_1517448501_1762 & f100;
   assign v3_1517448501_1822 = v3_1517448501_1819 & v3_1517448501_1820;
   assign v3_1517448501_1823 = ~v3_1517448501_1824;
   assign v3_1517448501_1824 = ~v3_1517448501_1767 & f101;
   assign v3_1517448501_1825 = v3_1517448501_1822 & v3_1517448501_1823;
   assign v3_1517448501_1826 = ~a_start_responder_0 & ~a_q;
   assign v3_1517448501_1827 = v3_1517448501_607 == v_kNb;
   assign v3_1517448501_1828 = v3_1517448501_1826 & v3_1517448501_1827;
   assign v3_1517448501_1829 = ~v3_1517448501_1830;
   assign v3_1517448501_1830 = f102 & ~v3_1517448501_1828;
   assign v3_1517448501_1831 = v3_1517448501_1825 & v3_1517448501_1829;
   assign v3_1517448501_1832 = ~a_start_responder_1 & ~a_q;
   assign v3_1517448501_1833 = v3_1517448501_1832 & v3_1517448501_1827;
   assign v3_1517448501_1834 = ~v3_1517448501_1835;
   assign v3_1517448501_1835 = f103 & ~v3_1517448501_1833;
   assign v3_1517448501_1836 = v3_1517448501_1831 & v3_1517448501_1834;
   assign v3_1517448501_1837 = ~a_start_responder_2 & ~a_q;
   assign v3_1517448501_1838 = v3_1517448501_1837 & v3_1517448501_1827;
   assign v3_1517448501_1839 = ~v3_1517448501_1840;
   assign v3_1517448501_1840 = f104 & ~v3_1517448501_1838;
   assign v3_1517448501_1841 = v3_1517448501_1836 & v3_1517448501_1839;
   assign v3_1517448501_1842 = ~v3_1517448501_1843;
   assign v3_1517448501_1843 = ~v3_1517448501_1828 & f105;
   assign v3_1517448501_1844 = v3_1517448501_1841 & v3_1517448501_1842;
   assign v3_1517448501_1845 = ~v3_1517448501_1846;
   assign v3_1517448501_1846 = ~v3_1517448501_1833 & f106;
   assign v3_1517448501_1847 = v3_1517448501_1844 & v3_1517448501_1845;
   assign v3_1517448501_1848 = ~v3_1517448501_1849;
   assign v3_1517448501_1849 = ~v3_1517448501_1838 & f107;
   assign v3_1517448501_1850 = v3_1517448501_1847 & v3_1517448501_1848;
   assign v3_1517448501_1851 = ~v3_1517448501_1852;
   assign v3_1517448501_1852 = ~v3_1517448501_1828 & f108;
   assign v3_1517448501_1853 = v3_1517448501_1850 & v3_1517448501_1851;
   assign v3_1517448501_1854 = ~v3_1517448501_1855;
   assign v3_1517448501_1855 = ~v3_1517448501_1833 & f109;
   assign v3_1517448501_1856 = v3_1517448501_1853 & v3_1517448501_1854;
   assign v3_1517448501_1857 = ~v3_1517448501_1858;
   assign v3_1517448501_1858 = ~v3_1517448501_1838 & f110;
   assign v3_1517448501_1859 = v3_1517448501_1856 & v3_1517448501_1857;
   assign v3_1517448501_1860 = a_wait_resp_initiator_0 & a_send_reply_responder_0;
   assign v3_1517448501_1861 = ~v3_1517448501_1862;
   assign v3_1517448501_1862 = f111 & ~v3_1517448501_1860;
   assign v3_1517448501_1863 = v3_1517448501_1859 & v3_1517448501_1861;
   assign v3_1517448501_1864 = a_wait_resp_initiator_1 & a_send_reply_responder_0;
   assign v3_1517448501_1865 = ~v3_1517448501_1866;
   assign v3_1517448501_1866 = f112 & ~v3_1517448501_1864;
   assign v3_1517448501_1867 = v3_1517448501_1863 & v3_1517448501_1865;
   assign v3_1517448501_1868 = a_wait_resp_initiator_2 & a_send_reply_responder_0;
   assign v3_1517448501_1869 = ~v3_1517448501_1870;
   assign v3_1517448501_1870 = f113 & ~v3_1517448501_1868;
   assign v3_1517448501_1871 = v3_1517448501_1867 & v3_1517448501_1869;
   assign v3_1517448501_1872 = a_send_reply_responder_0 & ~a_q;
   assign v3_1517448501_1873 = ~v3_1517448501_1874;
   assign v3_1517448501_1874 = f114 & ~v3_1517448501_1872;
   assign v3_1517448501_1875 = v3_1517448501_1871 & v3_1517448501_1873;
   assign v3_1517448501_1876 = a_wait_resp_initiator_0 & a_send_reply_responder_1;
   assign v3_1517448501_1877 = ~v3_1517448501_1878;
   assign v3_1517448501_1878 = f115 & ~v3_1517448501_1876;
   assign v3_1517448501_1879 = v3_1517448501_1875 & v3_1517448501_1877;
   assign v3_1517448501_1880 = a_wait_resp_initiator_1 & a_send_reply_responder_1;
   assign v3_1517448501_1881 = ~v3_1517448501_1882;
   assign v3_1517448501_1882 = f116 & ~v3_1517448501_1880;
   assign v3_1517448501_1883 = v3_1517448501_1879 & v3_1517448501_1881;
   assign v3_1517448501_1884 = a_wait_resp_initiator_2 & a_send_reply_responder_1;
   assign v3_1517448501_1885 = ~v3_1517448501_1886;
   assign v3_1517448501_1886 = f117 & ~v3_1517448501_1884;
   assign v3_1517448501_1887 = v3_1517448501_1883 & v3_1517448501_1885;
   assign v3_1517448501_1888 = a_send_reply_responder_1 & ~a_q;
   assign v3_1517448501_1889 = ~v3_1517448501_1890;
   assign v3_1517448501_1890 = f118 & ~v3_1517448501_1888;
   assign v3_1517448501_1891 = v3_1517448501_1887 & v3_1517448501_1889;
   assign v3_1517448501_1892 = a_wait_resp_initiator_0 & a_send_reply_responder_2;
   assign v3_1517448501_1893 = ~v3_1517448501_1894;
   assign v3_1517448501_1894 = f119 & ~v3_1517448501_1892;
   assign v3_1517448501_1895 = v3_1517448501_1891 & v3_1517448501_1893;
   assign v3_1517448501_1896 = a_wait_resp_initiator_1 & a_send_reply_responder_2;
   assign v3_1517448501_1897 = ~v3_1517448501_1898;
   assign v3_1517448501_1898 = f120 & ~v3_1517448501_1896;
   assign v3_1517448501_1899 = v3_1517448501_1895 & v3_1517448501_1897;
   assign v3_1517448501_1900 = a_wait_resp_initiator_2 & a_send_reply_responder_2;
   assign v3_1517448501_1901 = ~v3_1517448501_1902;
   assign v3_1517448501_1902 = f121 & ~v3_1517448501_1900;
   assign v3_1517448501_1903 = v3_1517448501_1899 & v3_1517448501_1901;
   assign v3_1517448501_1904 = a_send_reply_responder_2 & ~a_q;
   assign v3_1517448501_1905 = ~v3_1517448501_1906;
   assign v3_1517448501_1906 = f122 & ~v3_1517448501_1904;
   assign v3_1517448501_1907 = v3_1517448501_1903 & v3_1517448501_1905;
   assign v3_1517448501_1908 = a_wait_resp_initiator_0 & ~a_q;
   assign v3_1517448501_1909 = v3_1517448501_1908 & v3_1517448501_1756;
   assign v3_1517448501_1910 = ~v3_1517448501_1911;
   assign v3_1517448501_1911 = f123 & ~v3_1517448501_1909;
   assign v3_1517448501_1912 = v3_1517448501_1907 & v3_1517448501_1910;
   assign v3_1517448501_1913 = a_wait_resp_initiator_1 & ~a_q;
   assign v3_1517448501_1914 = v3_1517448501_1913 & v3_1517448501_1756;
   assign v3_1517448501_1915 = ~v3_1517448501_1916;
   assign v3_1517448501_1916 = f124 & ~v3_1517448501_1914;
   assign v3_1517448501_1917 = v3_1517448501_1912 & v3_1517448501_1915;
   assign v3_1517448501_1918 = a_wait_resp_initiator_2 & ~a_q;
   assign v3_1517448501_1919 = v3_1517448501_1918 & v3_1517448501_1756;
   assign v3_1517448501_1920 = ~v3_1517448501_1921;
   assign v3_1517448501_1921 = f125 & ~v3_1517448501_1919;
   assign v3_1517448501_1922 = v3_1517448501_1917 & v3_1517448501_1920;
   assign v3_1517448501_1923 = a_wait_resp_initiator_0 & ~a_q;
   assign v3_1517448501_1924 = v3_1517448501_1756 & v3_1517448501_1827;
   assign v3_1517448501_1925 = v3_1517448501_607 == v_k_Na_Nb__A;
   assign v3_1517448501_1926 = ~v3_1517448501_1927;
   assign v3_1517448501_1927 = ~v3_1517448501_1924 & ~v3_1517448501_1925;
   assign v3_1517448501_1928 = v3_1517448501_1923 & v3_1517448501_1926;
   assign v3_1517448501_1929 = ~v3_1517448501_1930;
   assign v3_1517448501_1930 = f126 & ~v3_1517448501_1928;
   assign v3_1517448501_1931 = v3_1517448501_1922 & v3_1517448501_1929;
   assign v3_1517448501_1932 = a_wait_resp_initiator_1 & ~a_q;
   assign v3_1517448501_1933 = v3_1517448501_1932 & v3_1517448501_1926;
   assign v3_1517448501_1934 = ~v3_1517448501_1935;
   assign v3_1517448501_1935 = f127 & ~v3_1517448501_1933;
   assign v3_1517448501_1936 = v3_1517448501_1931 & v3_1517448501_1934;
   assign v3_1517448501_1937 = a_wait_resp_initiator_2 & ~a_q;
   assign v3_1517448501_1938 = v3_1517448501_1937 & v3_1517448501_1926;
   assign v3_1517448501_1939 = ~v3_1517448501_1940;
   assign v3_1517448501_1940 = f128 & ~v3_1517448501_1938;
   assign v3_1517448501_1941 = v3_1517448501_1936 & v3_1517448501_1939;
   assign v3_1517448501_1942 = ~v3_1517448501_1943;
   assign v3_1517448501_1943 = ~v3_1517448501_1909 & f129;
   assign v3_1517448501_1944 = v3_1517448501_1941 & v3_1517448501_1942;
   assign v3_1517448501_1945 = ~v3_1517448501_1946;
   assign v3_1517448501_1946 = ~v3_1517448501_1914 & f130;
   assign v3_1517448501_1947 = v3_1517448501_1944 & v3_1517448501_1945;
   assign v3_1517448501_1948 = ~v3_1517448501_1949;
   assign v3_1517448501_1949 = ~v3_1517448501_1919 & f131;
   assign v3_1517448501_1950 = v3_1517448501_1947 & v3_1517448501_1948;
   assign v3_1517448501_1951 = a_commited_initiator_0 & a_wait_resp_responder_0;
   assign v3_1517448501_1952 = ~v3_1517448501_1953;
   assign v3_1517448501_1953 = f132 & ~v3_1517448501_1951;
   assign v3_1517448501_1954 = v3_1517448501_1950 & v3_1517448501_1952;
   assign v3_1517448501_1955 = a_commited_initiator_0 & a_wait_resp_responder_1;
   assign v3_1517448501_1956 = ~v3_1517448501_1957;
   assign v3_1517448501_1957 = f133 & ~v3_1517448501_1955;
   assign v3_1517448501_1958 = v3_1517448501_1954 & v3_1517448501_1956;
   assign v3_1517448501_1959 = a_commited_initiator_0 & a_wait_resp_responder_2;
   assign v3_1517448501_1960 = ~v3_1517448501_1961;
   assign v3_1517448501_1961 = f134 & ~v3_1517448501_1959;
   assign v3_1517448501_1962 = v3_1517448501_1958 & v3_1517448501_1960;
   assign v3_1517448501_1963 = a_commited_initiator_0 & ~a_q;
   assign v3_1517448501_1964 = ~v3_1517448501_1965;
   assign v3_1517448501_1965 = f135 & ~v3_1517448501_1963;
   assign v3_1517448501_1966 = v3_1517448501_1962 & v3_1517448501_1964;
   assign v3_1517448501_1967 = a_commited_initiator_1 & a_wait_resp_responder_0;
   assign v3_1517448501_1968 = ~v3_1517448501_1969;
   assign v3_1517448501_1969 = f136 & ~v3_1517448501_1967;
   assign v3_1517448501_1970 = v3_1517448501_1966 & v3_1517448501_1968;
   assign v3_1517448501_1971 = a_commited_initiator_1 & a_wait_resp_responder_1;
   assign v3_1517448501_1972 = ~v3_1517448501_1973;
   assign v3_1517448501_1973 = f137 & ~v3_1517448501_1971;
   assign v3_1517448501_1974 = v3_1517448501_1970 & v3_1517448501_1972;
   assign v3_1517448501_1975 = a_commited_initiator_1 & a_wait_resp_responder_2;
   assign v3_1517448501_1976 = ~v3_1517448501_1977;
   assign v3_1517448501_1977 = f138 & ~v3_1517448501_1975;
   assign v3_1517448501_1978 = v3_1517448501_1974 & v3_1517448501_1976;
   assign v3_1517448501_1979 = a_commited_initiator_1 & ~a_q;
   assign v3_1517448501_1980 = ~v3_1517448501_1981;
   assign v3_1517448501_1981 = f139 & ~v3_1517448501_1979;
   assign v3_1517448501_1982 = v3_1517448501_1978 & v3_1517448501_1980;
   assign v3_1517448501_1983 = a_commited_initiator_2 & a_wait_resp_responder_0;
   assign v3_1517448501_1984 = ~v3_1517448501_1985;
   assign v3_1517448501_1985 = f140 & ~v3_1517448501_1983;
   assign v3_1517448501_1986 = v3_1517448501_1982 & v3_1517448501_1984;
   assign v3_1517448501_1987 = a_commited_initiator_2 & a_wait_resp_responder_1;
   assign v3_1517448501_1988 = ~v3_1517448501_1989;
   assign v3_1517448501_1989 = f141 & ~v3_1517448501_1987;
   assign v3_1517448501_1990 = v3_1517448501_1986 & v3_1517448501_1988;
   assign v3_1517448501_1991 = a_commited_initiator_2 & a_wait_resp_responder_2;
   assign v3_1517448501_1992 = ~v3_1517448501_1993;
   assign v3_1517448501_1993 = f142 & ~v3_1517448501_1991;
   assign v3_1517448501_1994 = v3_1517448501_1990 & v3_1517448501_1992;
   assign v3_1517448501_1995 = a_commited_initiator_2 & ~a_q;
   assign v3_1517448501_1996 = ~v3_1517448501_1997;
   assign v3_1517448501_1997 = f143 & ~v3_1517448501_1995;
   assign v3_1517448501_1998 = v3_1517448501_1994 & v3_1517448501_1996;
   assign v3_1517448501_1999 = a_wait_resp_responder_0 & ~a_q;
   assign v3_1517448501_2000 = v3_1517448501_607 == v_k_Nb__B;
   assign v3_1517448501_2001 = ~v3_1517448501_2002;
   assign v3_1517448501_2002 = ~v3_1517448501_1827 & ~v3_1517448501_2000;
   assign v3_1517448501_2003 = v3_1517448501_1999 & v3_1517448501_2001;
   assign v3_1517448501_2004 = ~v3_1517448501_2005;
   assign v3_1517448501_2005 = f144 & ~v3_1517448501_2003;
   assign v3_1517448501_2006 = v3_1517448501_1998 & v3_1517448501_2004;
   assign v3_1517448501_2007 = a_wait_resp_responder_1 & ~a_q;
   assign v3_1517448501_2008 = v3_1517448501_2007 & v3_1517448501_2001;
   assign v3_1517448501_2009 = ~v3_1517448501_2010;
   assign v3_1517448501_2010 = f145 & ~v3_1517448501_2008;
   assign v3_1517448501_2011 = v3_1517448501_2006 & v3_1517448501_2009;
   assign v3_1517448501_2012 = a_wait_resp_responder_2 & ~a_q;
   assign v3_1517448501_2013 = v3_1517448501_2012 & v3_1517448501_2001;
   assign v3_1517448501_2014 = ~v3_1517448501_2015;
   assign v3_1517448501_2015 = f146 & ~v3_1517448501_2013;
   assign v3_1517448501_2016 = v3_1517448501_2011 & v3_1517448501_2014;
   assign v3_1517448501_2017 = ~v3_1517448501_2018;
   assign v3_1517448501_2018 = ~f000 & ~f001;
   assign v3_1517448501_2019 = ~v3_1517448501_2020;
   assign v3_1517448501_2020 = ~f002 & ~v3_1517448501_2017;
   assign v3_1517448501_2021 = ~v3_1517448501_2022;
   assign v3_1517448501_2022 = ~f003 & ~v3_1517448501_2019;
   assign v3_1517448501_2023 = ~v3_1517448501_2024;
   assign v3_1517448501_2024 = ~f004 & ~v3_1517448501_2021;
   assign v3_1517448501_2025 = ~v3_1517448501_2026;
   assign v3_1517448501_2026 = ~f005 & ~v3_1517448501_2023;
   assign v3_1517448501_2027 = ~v3_1517448501_2028;
   assign v3_1517448501_2028 = ~f006 & ~v3_1517448501_2025;
   assign v3_1517448501_2029 = ~v3_1517448501_2030;
   assign v3_1517448501_2030 = ~f007 & ~v3_1517448501_2027;
   assign v3_1517448501_2031 = ~v3_1517448501_2032;
   assign v3_1517448501_2032 = ~f008 & ~v3_1517448501_2029;
   assign v3_1517448501_2033 = ~v3_1517448501_2034;
   assign v3_1517448501_2034 = ~f009 & ~v3_1517448501_2031;
   assign v3_1517448501_2035 = ~v3_1517448501_2036;
   assign v3_1517448501_2036 = ~f010 & ~v3_1517448501_2033;
   assign v3_1517448501_2037 = ~v3_1517448501_2038;
   assign v3_1517448501_2038 = ~f011 & ~v3_1517448501_2035;
   assign v3_1517448501_2039 = ~v3_1517448501_2040;
   assign v3_1517448501_2040 = ~f012 & ~v3_1517448501_2037;
   assign v3_1517448501_2041 = ~v3_1517448501_2042;
   assign v3_1517448501_2042 = ~f013 & ~v3_1517448501_2039;
   assign v3_1517448501_2043 = ~v3_1517448501_2044;
   assign v3_1517448501_2044 = ~f014 & ~v3_1517448501_2041;
   assign v3_1517448501_2045 = ~v3_1517448501_2046;
   assign v3_1517448501_2046 = ~f015 & ~v3_1517448501_2043;
   assign v3_1517448501_2047 = ~v3_1517448501_2048;
   assign v3_1517448501_2048 = ~f016 & ~v3_1517448501_2045;
   assign v3_1517448501_2049 = ~v3_1517448501_2050;
   assign v3_1517448501_2050 = ~f017 & ~v3_1517448501_2047;
   assign v3_1517448501_2051 = ~v3_1517448501_2052;
   assign v3_1517448501_2052 = ~f018 & ~v3_1517448501_2049;
   assign v3_1517448501_2053 = ~v3_1517448501_2054;
   assign v3_1517448501_2054 = ~f019 & ~v3_1517448501_2051;
   assign v3_1517448501_2055 = ~v3_1517448501_2056;
   assign v3_1517448501_2056 = ~f020 & ~v3_1517448501_2053;
   assign v3_1517448501_2057 = ~v3_1517448501_2058;
   assign v3_1517448501_2058 = ~f021 & ~v3_1517448501_2055;
   assign v3_1517448501_2059 = ~v3_1517448501_2060;
   assign v3_1517448501_2060 = ~f022 & ~v3_1517448501_2057;
   assign v3_1517448501_2061 = ~v3_1517448501_2062;
   assign v3_1517448501_2062 = ~f023 & ~v3_1517448501_2059;
   assign v3_1517448501_2063 = ~v3_1517448501_2064;
   assign v3_1517448501_2064 = ~f024 & ~v3_1517448501_2061;
   assign v3_1517448501_2065 = ~v3_1517448501_2066;
   assign v3_1517448501_2066 = ~f025 & ~v3_1517448501_2063;
   assign v3_1517448501_2067 = ~v3_1517448501_2068;
   assign v3_1517448501_2068 = ~f026 & ~v3_1517448501_2065;
   assign v3_1517448501_2069 = ~v3_1517448501_2070;
   assign v3_1517448501_2070 = ~f027 & ~v3_1517448501_2067;
   assign v3_1517448501_2071 = ~v3_1517448501_2072;
   assign v3_1517448501_2072 = ~f028 & ~v3_1517448501_2069;
   assign v3_1517448501_2073 = ~v3_1517448501_2074;
   assign v3_1517448501_2074 = ~f029 & ~v3_1517448501_2071;
   assign v3_1517448501_2075 = ~v3_1517448501_2076;
   assign v3_1517448501_2076 = ~f030 & ~v3_1517448501_2073;
   assign v3_1517448501_2077 = ~v3_1517448501_2078;
   assign v3_1517448501_2078 = ~f031 & ~v3_1517448501_2075;
   assign v3_1517448501_2079 = ~v3_1517448501_2080;
   assign v3_1517448501_2080 = ~f032 & ~v3_1517448501_2077;
   assign v3_1517448501_2081 = ~v3_1517448501_2082;
   assign v3_1517448501_2082 = ~f033 & ~v3_1517448501_2079;
   assign v3_1517448501_2083 = ~v3_1517448501_2084;
   assign v3_1517448501_2084 = ~f034 & ~v3_1517448501_2081;
   assign v3_1517448501_2085 = ~v3_1517448501_2086;
   assign v3_1517448501_2086 = ~f035 & ~v3_1517448501_2083;
   assign v3_1517448501_2087 = ~v3_1517448501_2088;
   assign v3_1517448501_2088 = ~f036 & ~v3_1517448501_2085;
   assign v3_1517448501_2089 = ~v3_1517448501_2090;
   assign v3_1517448501_2090 = ~f037 & ~v3_1517448501_2087;
   assign v3_1517448501_2091 = ~v3_1517448501_2092;
   assign v3_1517448501_2092 = ~f038 & ~v3_1517448501_2089;
   assign v3_1517448501_2093 = ~v3_1517448501_2094;
   assign v3_1517448501_2094 = ~f039 & ~v3_1517448501_2091;
   assign v3_1517448501_2095 = ~v3_1517448501_2096;
   assign v3_1517448501_2096 = ~f040 & ~v3_1517448501_2093;
   assign v3_1517448501_2097 = ~v3_1517448501_2098;
   assign v3_1517448501_2098 = ~f041 & ~v3_1517448501_2095;
   assign v3_1517448501_2099 = ~v3_1517448501_2100;
   assign v3_1517448501_2100 = ~f042 & ~v3_1517448501_2097;
   assign v3_1517448501_2101 = ~v3_1517448501_2102;
   assign v3_1517448501_2102 = ~f043 & ~v3_1517448501_2099;
   assign v3_1517448501_2103 = ~v3_1517448501_2104;
   assign v3_1517448501_2104 = ~f044 & ~v3_1517448501_2101;
   assign v3_1517448501_2105 = ~v3_1517448501_2106;
   assign v3_1517448501_2106 = ~f045 & ~v3_1517448501_2103;
   assign v3_1517448501_2107 = ~v3_1517448501_2108;
   assign v3_1517448501_2108 = ~f046 & ~v3_1517448501_2105;
   assign v3_1517448501_2109 = ~v3_1517448501_2110;
   assign v3_1517448501_2110 = ~f047 & ~v3_1517448501_2107;
   assign v3_1517448501_2111 = ~v3_1517448501_2112;
   assign v3_1517448501_2112 = ~f048 & ~v3_1517448501_2109;
   assign v3_1517448501_2113 = ~v3_1517448501_2114;
   assign v3_1517448501_2114 = ~f049 & ~v3_1517448501_2111;
   assign v3_1517448501_2115 = ~v3_1517448501_2116;
   assign v3_1517448501_2116 = ~f050 & ~v3_1517448501_2113;
   assign v3_1517448501_2117 = ~v3_1517448501_2118;
   assign v3_1517448501_2118 = ~f051 & ~v3_1517448501_2115;
   assign v3_1517448501_2119 = ~v3_1517448501_2120;
   assign v3_1517448501_2120 = ~f052 & ~v3_1517448501_2117;
   assign v3_1517448501_2121 = ~v3_1517448501_2122;
   assign v3_1517448501_2122 = ~f053 & ~v3_1517448501_2119;
   assign v3_1517448501_2123 = ~v3_1517448501_2124;
   assign v3_1517448501_2124 = ~f054 & ~v3_1517448501_2121;
   assign v3_1517448501_2125 = ~v3_1517448501_2126;
   assign v3_1517448501_2126 = ~f055 & ~v3_1517448501_2123;
   assign v3_1517448501_2127 = ~v3_1517448501_2128;
   assign v3_1517448501_2128 = ~f056 & ~v3_1517448501_2125;
   assign v3_1517448501_2129 = ~v3_1517448501_2130;
   assign v3_1517448501_2130 = ~f057 & ~v3_1517448501_2127;
   assign v3_1517448501_2131 = ~v3_1517448501_2132;
   assign v3_1517448501_2132 = ~f058 & ~v3_1517448501_2129;
   assign v3_1517448501_2133 = ~v3_1517448501_2134;
   assign v3_1517448501_2134 = ~f059 & ~v3_1517448501_2131;
   assign v3_1517448501_2135 = ~v3_1517448501_2136;
   assign v3_1517448501_2136 = ~f060 & ~v3_1517448501_2133;
   assign v3_1517448501_2137 = ~v3_1517448501_2138;
   assign v3_1517448501_2138 = ~f061 & ~v3_1517448501_2135;
   assign v3_1517448501_2139 = ~v3_1517448501_2140;
   assign v3_1517448501_2140 = ~f062 & ~v3_1517448501_2137;
   assign v3_1517448501_2141 = ~v3_1517448501_2142;
   assign v3_1517448501_2142 = ~f063 & ~v3_1517448501_2139;
   assign v3_1517448501_2143 = ~v3_1517448501_2144;
   assign v3_1517448501_2144 = ~f064 & ~v3_1517448501_2141;
   assign v3_1517448501_2145 = ~v3_1517448501_2146;
   assign v3_1517448501_2146 = ~f065 & ~v3_1517448501_2143;
   assign v3_1517448501_2147 = ~v3_1517448501_2148;
   assign v3_1517448501_2148 = ~f066 & ~v3_1517448501_2145;
   assign v3_1517448501_2149 = ~v3_1517448501_2150;
   assign v3_1517448501_2150 = ~f067 & ~v3_1517448501_2147;
   assign v3_1517448501_2151 = ~v3_1517448501_2152;
   assign v3_1517448501_2152 = ~f068 & ~v3_1517448501_2149;
   assign v3_1517448501_2153 = ~v3_1517448501_2154;
   assign v3_1517448501_2154 = ~f069 & ~v3_1517448501_2151;
   assign v3_1517448501_2155 = ~v3_1517448501_2156;
   assign v3_1517448501_2156 = ~f070 & ~v3_1517448501_2153;
   assign v3_1517448501_2157 = ~v3_1517448501_2158;
   assign v3_1517448501_2158 = ~f071 & ~v3_1517448501_2155;
   assign v3_1517448501_2159 = ~v3_1517448501_2160;
   assign v3_1517448501_2160 = ~f072 & ~v3_1517448501_2157;
   assign v3_1517448501_2161 = ~v3_1517448501_2162;
   assign v3_1517448501_2162 = ~f073 & ~v3_1517448501_2159;
   assign v3_1517448501_2163 = ~v3_1517448501_2164;
   assign v3_1517448501_2164 = ~f074 & ~v3_1517448501_2161;
   assign v3_1517448501_2165 = ~v3_1517448501_2166;
   assign v3_1517448501_2166 = ~f075 & ~v3_1517448501_2163;
   assign v3_1517448501_2167 = ~v3_1517448501_2168;
   assign v3_1517448501_2168 = ~f076 & ~v3_1517448501_2165;
   assign v3_1517448501_2169 = ~v3_1517448501_2170;
   assign v3_1517448501_2170 = ~f077 & ~v3_1517448501_2167;
   assign v3_1517448501_2171 = ~v3_1517448501_2172;
   assign v3_1517448501_2172 = ~f078 & ~v3_1517448501_2169;
   assign v3_1517448501_2173 = ~v3_1517448501_2174;
   assign v3_1517448501_2174 = ~f079 & ~v3_1517448501_2171;
   assign v3_1517448501_2175 = ~v3_1517448501_2176;
   assign v3_1517448501_2176 = ~f080 & ~v3_1517448501_2173;
   assign v3_1517448501_2177 = ~v3_1517448501_2178;
   assign v3_1517448501_2178 = ~f081 & ~v3_1517448501_2175;
   assign v3_1517448501_2179 = ~v3_1517448501_2180;
   assign v3_1517448501_2180 = ~f082 & ~v3_1517448501_2177;
   assign v3_1517448501_2181 = ~v3_1517448501_2182;
   assign v3_1517448501_2182 = ~f083 & ~v3_1517448501_2179;
   assign v3_1517448501_2183 = ~v3_1517448501_2184;
   assign v3_1517448501_2184 = ~f084 & ~v3_1517448501_2181;
   assign v3_1517448501_2185 = ~v3_1517448501_2186;
   assign v3_1517448501_2186 = ~f085 & ~v3_1517448501_2183;
   assign v3_1517448501_2187 = ~v3_1517448501_2188;
   assign v3_1517448501_2188 = ~f086 & ~v3_1517448501_2185;
   assign v3_1517448501_2189 = ~v3_1517448501_2190;
   assign v3_1517448501_2190 = ~f087 & ~v3_1517448501_2187;
   assign v3_1517448501_2191 = ~v3_1517448501_2192;
   assign v3_1517448501_2192 = ~f088 & ~v3_1517448501_2189;
   assign v3_1517448501_2193 = ~v3_1517448501_2194;
   assign v3_1517448501_2194 = ~f089 & ~v3_1517448501_2191;
   assign v3_1517448501_2195 = ~v3_1517448501_2196;
   assign v3_1517448501_2196 = ~f090 & ~v3_1517448501_2193;
   assign v3_1517448501_2197 = ~v3_1517448501_2198;
   assign v3_1517448501_2198 = ~f091 & ~v3_1517448501_2195;
   assign v3_1517448501_2199 = ~v3_1517448501_2200;
   assign v3_1517448501_2200 = ~f092 & ~v3_1517448501_2197;
   assign v3_1517448501_2201 = ~v3_1517448501_2202;
   assign v3_1517448501_2202 = ~f093 & ~v3_1517448501_2199;
   assign v3_1517448501_2203 = ~v3_1517448501_2204;
   assign v3_1517448501_2204 = ~f094 & ~v3_1517448501_2201;
   assign v3_1517448501_2205 = ~v3_1517448501_2206;
   assign v3_1517448501_2206 = ~f095 & ~v3_1517448501_2203;
   assign v3_1517448501_2207 = ~v3_1517448501_2208;
   assign v3_1517448501_2208 = ~f096 & ~v3_1517448501_2205;
   assign v3_1517448501_2209 = ~v3_1517448501_2210;
   assign v3_1517448501_2210 = ~f097 & ~v3_1517448501_2207;
   assign v3_1517448501_2211 = ~v3_1517448501_2212;
   assign v3_1517448501_2212 = ~f098 & ~v3_1517448501_2209;
   assign v3_1517448501_2213 = ~v3_1517448501_2214;
   assign v3_1517448501_2214 = ~f099 & ~v3_1517448501_2211;
   assign v3_1517448501_2215 = ~v3_1517448501_2216;
   assign v3_1517448501_2216 = ~f100 & ~v3_1517448501_2213;
   assign v3_1517448501_2217 = ~v3_1517448501_2218;
   assign v3_1517448501_2218 = ~f101 & ~v3_1517448501_2215;
   assign v3_1517448501_2219 = ~v3_1517448501_2220;
   assign v3_1517448501_2220 = ~f102 & ~v3_1517448501_2217;
   assign v3_1517448501_2221 = ~v3_1517448501_2222;
   assign v3_1517448501_2222 = ~f103 & ~v3_1517448501_2219;
   assign v3_1517448501_2223 = ~v3_1517448501_2224;
   assign v3_1517448501_2224 = ~f104 & ~v3_1517448501_2221;
   assign v3_1517448501_2225 = ~v3_1517448501_2226;
   assign v3_1517448501_2226 = ~f105 & ~v3_1517448501_2223;
   assign v3_1517448501_2227 = ~v3_1517448501_2228;
   assign v3_1517448501_2228 = ~f106 & ~v3_1517448501_2225;
   assign v3_1517448501_2229 = ~v3_1517448501_2230;
   assign v3_1517448501_2230 = ~f107 & ~v3_1517448501_2227;
   assign v3_1517448501_2231 = ~v3_1517448501_2232;
   assign v3_1517448501_2232 = ~f108 & ~v3_1517448501_2229;
   assign v3_1517448501_2233 = ~v3_1517448501_2234;
   assign v3_1517448501_2234 = ~f109 & ~v3_1517448501_2231;
   assign v3_1517448501_2235 = ~v3_1517448501_2236;
   assign v3_1517448501_2236 = ~f110 & ~v3_1517448501_2233;
   assign v3_1517448501_2237 = ~v3_1517448501_2238;
   assign v3_1517448501_2238 = ~f111 & ~v3_1517448501_2235;
   assign v3_1517448501_2239 = ~v3_1517448501_2240;
   assign v3_1517448501_2240 = ~f112 & ~v3_1517448501_2237;
   assign v3_1517448501_2241 = ~v3_1517448501_2242;
   assign v3_1517448501_2242 = ~f113 & ~v3_1517448501_2239;
   assign v3_1517448501_2243 = ~v3_1517448501_2244;
   assign v3_1517448501_2244 = ~f114 & ~v3_1517448501_2241;
   assign v3_1517448501_2245 = ~v3_1517448501_2246;
   assign v3_1517448501_2246 = ~f115 & ~v3_1517448501_2243;
   assign v3_1517448501_2247 = ~v3_1517448501_2248;
   assign v3_1517448501_2248 = ~f116 & ~v3_1517448501_2245;
   assign v3_1517448501_2249 = ~v3_1517448501_2250;
   assign v3_1517448501_2250 = ~f117 & ~v3_1517448501_2247;
   assign v3_1517448501_2251 = ~v3_1517448501_2252;
   assign v3_1517448501_2252 = ~f118 & ~v3_1517448501_2249;
   assign v3_1517448501_2253 = ~v3_1517448501_2254;
   assign v3_1517448501_2254 = ~f119 & ~v3_1517448501_2251;
   assign v3_1517448501_2255 = ~v3_1517448501_2256;
   assign v3_1517448501_2256 = ~f120 & ~v3_1517448501_2253;
   assign v3_1517448501_2257 = ~v3_1517448501_2258;
   assign v3_1517448501_2258 = ~f121 & ~v3_1517448501_2255;
   assign v3_1517448501_2259 = ~v3_1517448501_2260;
   assign v3_1517448501_2260 = ~f122 & ~v3_1517448501_2257;
   assign v3_1517448501_2261 = ~v3_1517448501_2262;
   assign v3_1517448501_2262 = ~f123 & ~v3_1517448501_2259;
   assign v3_1517448501_2263 = ~v3_1517448501_2264;
   assign v3_1517448501_2264 = ~f124 & ~v3_1517448501_2261;
   assign v3_1517448501_2265 = ~v3_1517448501_2266;
   assign v3_1517448501_2266 = ~f125 & ~v3_1517448501_2263;
   assign v3_1517448501_2267 = ~v3_1517448501_2268;
   assign v3_1517448501_2268 = ~f126 & ~v3_1517448501_2265;
   assign v3_1517448501_2269 = ~v3_1517448501_2270;
   assign v3_1517448501_2270 = ~f127 & ~v3_1517448501_2267;
   assign v3_1517448501_2271 = ~v3_1517448501_2272;
   assign v3_1517448501_2272 = ~f128 & ~v3_1517448501_2269;
   assign v3_1517448501_2273 = ~v3_1517448501_2274;
   assign v3_1517448501_2274 = ~f129 & ~v3_1517448501_2271;
   assign v3_1517448501_2275 = ~v3_1517448501_2276;
   assign v3_1517448501_2276 = ~f130 & ~v3_1517448501_2273;
   assign v3_1517448501_2277 = ~v3_1517448501_2278;
   assign v3_1517448501_2278 = ~f131 & ~v3_1517448501_2275;
   assign v3_1517448501_2279 = ~v3_1517448501_2280;
   assign v3_1517448501_2280 = ~f132 & ~v3_1517448501_2277;
   assign v3_1517448501_2281 = ~v3_1517448501_2282;
   assign v3_1517448501_2282 = ~f133 & ~v3_1517448501_2279;
   assign v3_1517448501_2283 = ~v3_1517448501_2284;
   assign v3_1517448501_2284 = ~f134 & ~v3_1517448501_2281;
   assign v3_1517448501_2285 = ~v3_1517448501_2286;
   assign v3_1517448501_2286 = ~f135 & ~v3_1517448501_2283;
   assign v3_1517448501_2287 = ~v3_1517448501_2288;
   assign v3_1517448501_2288 = ~f136 & ~v3_1517448501_2285;
   assign v3_1517448501_2289 = ~v3_1517448501_2290;
   assign v3_1517448501_2290 = ~f137 & ~v3_1517448501_2287;
   assign v3_1517448501_2291 = ~v3_1517448501_2292;
   assign v3_1517448501_2292 = ~f138 & ~v3_1517448501_2289;
   assign v3_1517448501_2293 = ~v3_1517448501_2294;
   assign v3_1517448501_2294 = ~f139 & ~v3_1517448501_2291;
   assign v3_1517448501_2295 = ~v3_1517448501_2296;
   assign v3_1517448501_2296 = ~f140 & ~v3_1517448501_2293;
   assign v3_1517448501_2297 = ~v3_1517448501_2298;
   assign v3_1517448501_2298 = ~f141 & ~v3_1517448501_2295;
   assign v3_1517448501_2299 = ~v3_1517448501_2300;
   assign v3_1517448501_2300 = ~f142 & ~v3_1517448501_2297;
   assign v3_1517448501_2301 = ~v3_1517448501_2302;
   assign v3_1517448501_2302 = ~f143 & ~v3_1517448501_2299;
   assign v3_1517448501_2303 = ~v3_1517448501_2304;
   assign v3_1517448501_2304 = ~f144 & ~v3_1517448501_2301;
   assign v3_1517448501_2305 = ~v3_1517448501_2306;
   assign v3_1517448501_2306 = ~f145 & ~v3_1517448501_2303;
   assign v3_1517448501_2307 = ~v3_1517448501_2308;
   assign v3_1517448501_2308 = ~f146 & ~v3_1517448501_2305;
   assign v3_1517448501_2309 = v3_1517448501_2016 & v3_1517448501_2307;
   assign v3_1517448501_2310 = f000 & f001;
   assign v3_1517448501_2311 = f002 & v3_1517448501_2017;
   assign v3_1517448501_2312 = ~v3_1517448501_2313;
   assign v3_1517448501_2313 = ~v3_1517448501_2310 & ~v3_1517448501_2311;
   assign v3_1517448501_2314 = f003 & v3_1517448501_2019;
   assign v3_1517448501_2315 = ~v3_1517448501_2316;
   assign v3_1517448501_2316 = ~v3_1517448501_2312 & ~v3_1517448501_2314;
   assign v3_1517448501_2317 = f004 & v3_1517448501_2021;
   assign v3_1517448501_2318 = ~v3_1517448501_2319;
   assign v3_1517448501_2319 = ~v3_1517448501_2315 & ~v3_1517448501_2317;
   assign v3_1517448501_2320 = f005 & v3_1517448501_2023;
   assign v3_1517448501_2321 = ~v3_1517448501_2322;
   assign v3_1517448501_2322 = ~v3_1517448501_2318 & ~v3_1517448501_2320;
   assign v3_1517448501_2323 = f006 & v3_1517448501_2025;
   assign v3_1517448501_2324 = ~v3_1517448501_2325;
   assign v3_1517448501_2325 = ~v3_1517448501_2321 & ~v3_1517448501_2323;
   assign v3_1517448501_2326 = f007 & v3_1517448501_2027;
   assign v3_1517448501_2327 = ~v3_1517448501_2328;
   assign v3_1517448501_2328 = ~v3_1517448501_2324 & ~v3_1517448501_2326;
   assign v3_1517448501_2329 = f008 & v3_1517448501_2029;
   assign v3_1517448501_2330 = ~v3_1517448501_2331;
   assign v3_1517448501_2331 = ~v3_1517448501_2327 & ~v3_1517448501_2329;
   assign v3_1517448501_2332 = f009 & v3_1517448501_2031;
   assign v3_1517448501_2333 = ~v3_1517448501_2334;
   assign v3_1517448501_2334 = ~v3_1517448501_2330 & ~v3_1517448501_2332;
   assign v3_1517448501_2335 = f010 & v3_1517448501_2033;
   assign v3_1517448501_2336 = ~v3_1517448501_2337;
   assign v3_1517448501_2337 = ~v3_1517448501_2333 & ~v3_1517448501_2335;
   assign v3_1517448501_2338 = f011 & v3_1517448501_2035;
   assign v3_1517448501_2339 = ~v3_1517448501_2340;
   assign v3_1517448501_2340 = ~v3_1517448501_2336 & ~v3_1517448501_2338;
   assign v3_1517448501_2341 = f012 & v3_1517448501_2037;
   assign v3_1517448501_2342 = ~v3_1517448501_2343;
   assign v3_1517448501_2343 = ~v3_1517448501_2339 & ~v3_1517448501_2341;
   assign v3_1517448501_2344 = f013 & v3_1517448501_2039;
   assign v3_1517448501_2345 = ~v3_1517448501_2346;
   assign v3_1517448501_2346 = ~v3_1517448501_2342 & ~v3_1517448501_2344;
   assign v3_1517448501_2347 = f014 & v3_1517448501_2041;
   assign v3_1517448501_2348 = ~v3_1517448501_2349;
   assign v3_1517448501_2349 = ~v3_1517448501_2345 & ~v3_1517448501_2347;
   assign v3_1517448501_2350 = f015 & v3_1517448501_2043;
   assign v3_1517448501_2351 = ~v3_1517448501_2352;
   assign v3_1517448501_2352 = ~v3_1517448501_2348 & ~v3_1517448501_2350;
   assign v3_1517448501_2353 = f016 & v3_1517448501_2045;
   assign v3_1517448501_2354 = ~v3_1517448501_2355;
   assign v3_1517448501_2355 = ~v3_1517448501_2351 & ~v3_1517448501_2353;
   assign v3_1517448501_2356 = f017 & v3_1517448501_2047;
   assign v3_1517448501_2357 = ~v3_1517448501_2358;
   assign v3_1517448501_2358 = ~v3_1517448501_2354 & ~v3_1517448501_2356;
   assign v3_1517448501_2359 = f018 & v3_1517448501_2049;
   assign v3_1517448501_2360 = ~v3_1517448501_2361;
   assign v3_1517448501_2361 = ~v3_1517448501_2357 & ~v3_1517448501_2359;
   assign v3_1517448501_2362 = f019 & v3_1517448501_2051;
   assign v3_1517448501_2363 = ~v3_1517448501_2364;
   assign v3_1517448501_2364 = ~v3_1517448501_2360 & ~v3_1517448501_2362;
   assign v3_1517448501_2365 = f020 & v3_1517448501_2053;
   assign v3_1517448501_2366 = ~v3_1517448501_2367;
   assign v3_1517448501_2367 = ~v3_1517448501_2363 & ~v3_1517448501_2365;
   assign v3_1517448501_2368 = f021 & v3_1517448501_2055;
   assign v3_1517448501_2369 = ~v3_1517448501_2370;
   assign v3_1517448501_2370 = ~v3_1517448501_2366 & ~v3_1517448501_2368;
   assign v3_1517448501_2371 = f022 & v3_1517448501_2057;
   assign v3_1517448501_2372 = ~v3_1517448501_2373;
   assign v3_1517448501_2373 = ~v3_1517448501_2369 & ~v3_1517448501_2371;
   assign v3_1517448501_2374 = f023 & v3_1517448501_2059;
   assign v3_1517448501_2375 = ~v3_1517448501_2376;
   assign v3_1517448501_2376 = ~v3_1517448501_2372 & ~v3_1517448501_2374;
   assign v3_1517448501_2377 = f024 & v3_1517448501_2061;
   assign v3_1517448501_2378 = ~v3_1517448501_2379;
   assign v3_1517448501_2379 = ~v3_1517448501_2375 & ~v3_1517448501_2377;
   assign v3_1517448501_2380 = f025 & v3_1517448501_2063;
   assign v3_1517448501_2381 = ~v3_1517448501_2382;
   assign v3_1517448501_2382 = ~v3_1517448501_2378 & ~v3_1517448501_2380;
   assign v3_1517448501_2383 = f026 & v3_1517448501_2065;
   assign v3_1517448501_2384 = ~v3_1517448501_2385;
   assign v3_1517448501_2385 = ~v3_1517448501_2381 & ~v3_1517448501_2383;
   assign v3_1517448501_2386 = f027 & v3_1517448501_2067;
   assign v3_1517448501_2387 = ~v3_1517448501_2388;
   assign v3_1517448501_2388 = ~v3_1517448501_2384 & ~v3_1517448501_2386;
   assign v3_1517448501_2389 = f028 & v3_1517448501_2069;
   assign v3_1517448501_2390 = ~v3_1517448501_2391;
   assign v3_1517448501_2391 = ~v3_1517448501_2387 & ~v3_1517448501_2389;
   assign v3_1517448501_2392 = f029 & v3_1517448501_2071;
   assign v3_1517448501_2393 = ~v3_1517448501_2394;
   assign v3_1517448501_2394 = ~v3_1517448501_2390 & ~v3_1517448501_2392;
   assign v3_1517448501_2395 = f030 & v3_1517448501_2073;
   assign v3_1517448501_2396 = ~v3_1517448501_2397;
   assign v3_1517448501_2397 = ~v3_1517448501_2393 & ~v3_1517448501_2395;
   assign v3_1517448501_2398 = f031 & v3_1517448501_2075;
   assign v3_1517448501_2399 = ~v3_1517448501_2400;
   assign v3_1517448501_2400 = ~v3_1517448501_2396 & ~v3_1517448501_2398;
   assign v3_1517448501_2401 = f032 & v3_1517448501_2077;
   assign v3_1517448501_2402 = ~v3_1517448501_2403;
   assign v3_1517448501_2403 = ~v3_1517448501_2399 & ~v3_1517448501_2401;
   assign v3_1517448501_2404 = f033 & v3_1517448501_2079;
   assign v3_1517448501_2405 = ~v3_1517448501_2406;
   assign v3_1517448501_2406 = ~v3_1517448501_2402 & ~v3_1517448501_2404;
   assign v3_1517448501_2407 = f034 & v3_1517448501_2081;
   assign v3_1517448501_2408 = ~v3_1517448501_2409;
   assign v3_1517448501_2409 = ~v3_1517448501_2405 & ~v3_1517448501_2407;
   assign v3_1517448501_2410 = f035 & v3_1517448501_2083;
   assign v3_1517448501_2411 = ~v3_1517448501_2412;
   assign v3_1517448501_2412 = ~v3_1517448501_2408 & ~v3_1517448501_2410;
   assign v3_1517448501_2413 = f036 & v3_1517448501_2085;
   assign v3_1517448501_2414 = ~v3_1517448501_2415;
   assign v3_1517448501_2415 = ~v3_1517448501_2411 & ~v3_1517448501_2413;
   assign v3_1517448501_2416 = f037 & v3_1517448501_2087;
   assign v3_1517448501_2417 = ~v3_1517448501_2418;
   assign v3_1517448501_2418 = ~v3_1517448501_2414 & ~v3_1517448501_2416;
   assign v3_1517448501_2419 = f038 & v3_1517448501_2089;
   assign v3_1517448501_2420 = ~v3_1517448501_2421;
   assign v3_1517448501_2421 = ~v3_1517448501_2417 & ~v3_1517448501_2419;
   assign v3_1517448501_2422 = f039 & v3_1517448501_2091;
   assign v3_1517448501_2423 = ~v3_1517448501_2424;
   assign v3_1517448501_2424 = ~v3_1517448501_2420 & ~v3_1517448501_2422;
   assign v3_1517448501_2425 = f040 & v3_1517448501_2093;
   assign v3_1517448501_2426 = ~v3_1517448501_2427;
   assign v3_1517448501_2427 = ~v3_1517448501_2423 & ~v3_1517448501_2425;
   assign v3_1517448501_2428 = f041 & v3_1517448501_2095;
   assign v3_1517448501_2429 = ~v3_1517448501_2430;
   assign v3_1517448501_2430 = ~v3_1517448501_2426 & ~v3_1517448501_2428;
   assign v3_1517448501_2431 = f042 & v3_1517448501_2097;
   assign v3_1517448501_2432 = ~v3_1517448501_2433;
   assign v3_1517448501_2433 = ~v3_1517448501_2429 & ~v3_1517448501_2431;
   assign v3_1517448501_2434 = f043 & v3_1517448501_2099;
   assign v3_1517448501_2435 = ~v3_1517448501_2436;
   assign v3_1517448501_2436 = ~v3_1517448501_2432 & ~v3_1517448501_2434;
   assign v3_1517448501_2437 = f044 & v3_1517448501_2101;
   assign v3_1517448501_2438 = ~v3_1517448501_2439;
   assign v3_1517448501_2439 = ~v3_1517448501_2435 & ~v3_1517448501_2437;
   assign v3_1517448501_2440 = f045 & v3_1517448501_2103;
   assign v3_1517448501_2441 = ~v3_1517448501_2442;
   assign v3_1517448501_2442 = ~v3_1517448501_2438 & ~v3_1517448501_2440;
   assign v3_1517448501_2443 = f046 & v3_1517448501_2105;
   assign v3_1517448501_2444 = ~v3_1517448501_2445;
   assign v3_1517448501_2445 = ~v3_1517448501_2441 & ~v3_1517448501_2443;
   assign v3_1517448501_2446 = f047 & v3_1517448501_2107;
   assign v3_1517448501_2447 = ~v3_1517448501_2448;
   assign v3_1517448501_2448 = ~v3_1517448501_2444 & ~v3_1517448501_2446;
   assign v3_1517448501_2449 = f048 & v3_1517448501_2109;
   assign v3_1517448501_2450 = ~v3_1517448501_2451;
   assign v3_1517448501_2451 = ~v3_1517448501_2447 & ~v3_1517448501_2449;
   assign v3_1517448501_2452 = f049 & v3_1517448501_2111;
   assign v3_1517448501_2453 = ~v3_1517448501_2454;
   assign v3_1517448501_2454 = ~v3_1517448501_2450 & ~v3_1517448501_2452;
   assign v3_1517448501_2455 = f050 & v3_1517448501_2113;
   assign v3_1517448501_2456 = ~v3_1517448501_2457;
   assign v3_1517448501_2457 = ~v3_1517448501_2453 & ~v3_1517448501_2455;
   assign v3_1517448501_2458 = f051 & v3_1517448501_2115;
   assign v3_1517448501_2459 = ~v3_1517448501_2460;
   assign v3_1517448501_2460 = ~v3_1517448501_2456 & ~v3_1517448501_2458;
   assign v3_1517448501_2461 = f052 & v3_1517448501_2117;
   assign v3_1517448501_2462 = ~v3_1517448501_2463;
   assign v3_1517448501_2463 = ~v3_1517448501_2459 & ~v3_1517448501_2461;
   assign v3_1517448501_2464 = f053 & v3_1517448501_2119;
   assign v3_1517448501_2465 = ~v3_1517448501_2466;
   assign v3_1517448501_2466 = ~v3_1517448501_2462 & ~v3_1517448501_2464;
   assign v3_1517448501_2467 = f054 & v3_1517448501_2121;
   assign v3_1517448501_2468 = ~v3_1517448501_2469;
   assign v3_1517448501_2469 = ~v3_1517448501_2465 & ~v3_1517448501_2467;
   assign v3_1517448501_2470 = f055 & v3_1517448501_2123;
   assign v3_1517448501_2471 = ~v3_1517448501_2472;
   assign v3_1517448501_2472 = ~v3_1517448501_2468 & ~v3_1517448501_2470;
   assign v3_1517448501_2473 = f056 & v3_1517448501_2125;
   assign v3_1517448501_2474 = ~v3_1517448501_2475;
   assign v3_1517448501_2475 = ~v3_1517448501_2471 & ~v3_1517448501_2473;
   assign v3_1517448501_2476 = f057 & v3_1517448501_2127;
   assign v3_1517448501_2477 = ~v3_1517448501_2478;
   assign v3_1517448501_2478 = ~v3_1517448501_2474 & ~v3_1517448501_2476;
   assign v3_1517448501_2479 = f058 & v3_1517448501_2129;
   assign v3_1517448501_2480 = ~v3_1517448501_2481;
   assign v3_1517448501_2481 = ~v3_1517448501_2477 & ~v3_1517448501_2479;
   assign v3_1517448501_2482 = f059 & v3_1517448501_2131;
   assign v3_1517448501_2483 = ~v3_1517448501_2484;
   assign v3_1517448501_2484 = ~v3_1517448501_2480 & ~v3_1517448501_2482;
   assign v3_1517448501_2485 = f060 & v3_1517448501_2133;
   assign v3_1517448501_2486 = ~v3_1517448501_2487;
   assign v3_1517448501_2487 = ~v3_1517448501_2483 & ~v3_1517448501_2485;
   assign v3_1517448501_2488 = f061 & v3_1517448501_2135;
   assign v3_1517448501_2489 = ~v3_1517448501_2490;
   assign v3_1517448501_2490 = ~v3_1517448501_2486 & ~v3_1517448501_2488;
   assign v3_1517448501_2491 = f062 & v3_1517448501_2137;
   assign v3_1517448501_2492 = ~v3_1517448501_2493;
   assign v3_1517448501_2493 = ~v3_1517448501_2489 & ~v3_1517448501_2491;
   assign v3_1517448501_2494 = f063 & v3_1517448501_2139;
   assign v3_1517448501_2495 = ~v3_1517448501_2496;
   assign v3_1517448501_2496 = ~v3_1517448501_2492 & ~v3_1517448501_2494;
   assign v3_1517448501_2497 = f064 & v3_1517448501_2141;
   assign v3_1517448501_2498 = ~v3_1517448501_2499;
   assign v3_1517448501_2499 = ~v3_1517448501_2495 & ~v3_1517448501_2497;
   assign v3_1517448501_2500 = f065 & v3_1517448501_2143;
   assign v3_1517448501_2501 = ~v3_1517448501_2502;
   assign v3_1517448501_2502 = ~v3_1517448501_2498 & ~v3_1517448501_2500;
   assign v3_1517448501_2503 = f066 & v3_1517448501_2145;
   assign v3_1517448501_2504 = ~v3_1517448501_2505;
   assign v3_1517448501_2505 = ~v3_1517448501_2501 & ~v3_1517448501_2503;
   assign v3_1517448501_2506 = f067 & v3_1517448501_2147;
   assign v3_1517448501_2507 = ~v3_1517448501_2508;
   assign v3_1517448501_2508 = ~v3_1517448501_2504 & ~v3_1517448501_2506;
   assign v3_1517448501_2509 = f068 & v3_1517448501_2149;
   assign v3_1517448501_2510 = ~v3_1517448501_2511;
   assign v3_1517448501_2511 = ~v3_1517448501_2507 & ~v3_1517448501_2509;
   assign v3_1517448501_2512 = f069 & v3_1517448501_2151;
   assign v3_1517448501_2513 = ~v3_1517448501_2514;
   assign v3_1517448501_2514 = ~v3_1517448501_2510 & ~v3_1517448501_2512;
   assign v3_1517448501_2515 = f070 & v3_1517448501_2153;
   assign v3_1517448501_2516 = ~v3_1517448501_2517;
   assign v3_1517448501_2517 = ~v3_1517448501_2513 & ~v3_1517448501_2515;
   assign v3_1517448501_2518 = f071 & v3_1517448501_2155;
   assign v3_1517448501_2519 = ~v3_1517448501_2520;
   assign v3_1517448501_2520 = ~v3_1517448501_2516 & ~v3_1517448501_2518;
   assign v3_1517448501_2521 = f072 & v3_1517448501_2157;
   assign v3_1517448501_2522 = ~v3_1517448501_2523;
   assign v3_1517448501_2523 = ~v3_1517448501_2519 & ~v3_1517448501_2521;
   assign v3_1517448501_2524 = f073 & v3_1517448501_2159;
   assign v3_1517448501_2525 = ~v3_1517448501_2526;
   assign v3_1517448501_2526 = ~v3_1517448501_2522 & ~v3_1517448501_2524;
   assign v3_1517448501_2527 = f074 & v3_1517448501_2161;
   assign v3_1517448501_2528 = ~v3_1517448501_2529;
   assign v3_1517448501_2529 = ~v3_1517448501_2525 & ~v3_1517448501_2527;
   assign v3_1517448501_2530 = f075 & v3_1517448501_2163;
   assign v3_1517448501_2531 = ~v3_1517448501_2532;
   assign v3_1517448501_2532 = ~v3_1517448501_2528 & ~v3_1517448501_2530;
   assign v3_1517448501_2533 = f076 & v3_1517448501_2165;
   assign v3_1517448501_2534 = ~v3_1517448501_2535;
   assign v3_1517448501_2535 = ~v3_1517448501_2531 & ~v3_1517448501_2533;
   assign v3_1517448501_2536 = f077 & v3_1517448501_2167;
   assign v3_1517448501_2537 = ~v3_1517448501_2538;
   assign v3_1517448501_2538 = ~v3_1517448501_2534 & ~v3_1517448501_2536;
   assign v3_1517448501_2539 = f078 & v3_1517448501_2169;
   assign v3_1517448501_2540 = ~v3_1517448501_2541;
   assign v3_1517448501_2541 = ~v3_1517448501_2537 & ~v3_1517448501_2539;
   assign v3_1517448501_2542 = f079 & v3_1517448501_2171;
   assign v3_1517448501_2543 = ~v3_1517448501_2544;
   assign v3_1517448501_2544 = ~v3_1517448501_2540 & ~v3_1517448501_2542;
   assign v3_1517448501_2545 = f080 & v3_1517448501_2173;
   assign v3_1517448501_2546 = ~v3_1517448501_2547;
   assign v3_1517448501_2547 = ~v3_1517448501_2543 & ~v3_1517448501_2545;
   assign v3_1517448501_2548 = f081 & v3_1517448501_2175;
   assign v3_1517448501_2549 = ~v3_1517448501_2550;
   assign v3_1517448501_2550 = ~v3_1517448501_2546 & ~v3_1517448501_2548;
   assign v3_1517448501_2551 = f082 & v3_1517448501_2177;
   assign v3_1517448501_2552 = ~v3_1517448501_2553;
   assign v3_1517448501_2553 = ~v3_1517448501_2549 & ~v3_1517448501_2551;
   assign v3_1517448501_2554 = f083 & v3_1517448501_2179;
   assign v3_1517448501_2555 = ~v3_1517448501_2556;
   assign v3_1517448501_2556 = ~v3_1517448501_2552 & ~v3_1517448501_2554;
   assign v3_1517448501_2557 = f084 & v3_1517448501_2181;
   assign v3_1517448501_2558 = ~v3_1517448501_2559;
   assign v3_1517448501_2559 = ~v3_1517448501_2555 & ~v3_1517448501_2557;
   assign v3_1517448501_2560 = f085 & v3_1517448501_2183;
   assign v3_1517448501_2561 = ~v3_1517448501_2562;
   assign v3_1517448501_2562 = ~v3_1517448501_2558 & ~v3_1517448501_2560;
   assign v3_1517448501_2563 = f086 & v3_1517448501_2185;
   assign v3_1517448501_2564 = ~v3_1517448501_2565;
   assign v3_1517448501_2565 = ~v3_1517448501_2561 & ~v3_1517448501_2563;
   assign v3_1517448501_2566 = f087 & v3_1517448501_2187;
   assign v3_1517448501_2567 = ~v3_1517448501_2568;
   assign v3_1517448501_2568 = ~v3_1517448501_2564 & ~v3_1517448501_2566;
   assign v3_1517448501_2569 = f088 & v3_1517448501_2189;
   assign v3_1517448501_2570 = ~v3_1517448501_2571;
   assign v3_1517448501_2571 = ~v3_1517448501_2567 & ~v3_1517448501_2569;
   assign v3_1517448501_2572 = f089 & v3_1517448501_2191;
   assign v3_1517448501_2573 = ~v3_1517448501_2574;
   assign v3_1517448501_2574 = ~v3_1517448501_2570 & ~v3_1517448501_2572;
   assign v3_1517448501_2575 = f090 & v3_1517448501_2193;
   assign v3_1517448501_2576 = ~v3_1517448501_2577;
   assign v3_1517448501_2577 = ~v3_1517448501_2573 & ~v3_1517448501_2575;
   assign v3_1517448501_2578 = f091 & v3_1517448501_2195;
   assign v3_1517448501_2579 = ~v3_1517448501_2580;
   assign v3_1517448501_2580 = ~v3_1517448501_2576 & ~v3_1517448501_2578;
   assign v3_1517448501_2581 = f092 & v3_1517448501_2197;
   assign v3_1517448501_2582 = ~v3_1517448501_2583;
   assign v3_1517448501_2583 = ~v3_1517448501_2579 & ~v3_1517448501_2581;
   assign v3_1517448501_2584 = f093 & v3_1517448501_2199;
   assign v3_1517448501_2585 = ~v3_1517448501_2586;
   assign v3_1517448501_2586 = ~v3_1517448501_2582 & ~v3_1517448501_2584;
   assign v3_1517448501_2587 = f094 & v3_1517448501_2201;
   assign v3_1517448501_2588 = ~v3_1517448501_2589;
   assign v3_1517448501_2589 = ~v3_1517448501_2585 & ~v3_1517448501_2587;
   assign v3_1517448501_2590 = f095 & v3_1517448501_2203;
   assign v3_1517448501_2591 = ~v3_1517448501_2592;
   assign v3_1517448501_2592 = ~v3_1517448501_2588 & ~v3_1517448501_2590;
   assign v3_1517448501_2593 = f096 & v3_1517448501_2205;
   assign v3_1517448501_2594 = ~v3_1517448501_2595;
   assign v3_1517448501_2595 = ~v3_1517448501_2591 & ~v3_1517448501_2593;
   assign v3_1517448501_2596 = f097 & v3_1517448501_2207;
   assign v3_1517448501_2597 = ~v3_1517448501_2598;
   assign v3_1517448501_2598 = ~v3_1517448501_2594 & ~v3_1517448501_2596;
   assign v3_1517448501_2599 = f098 & v3_1517448501_2209;
   assign v3_1517448501_2600 = ~v3_1517448501_2601;
   assign v3_1517448501_2601 = ~v3_1517448501_2597 & ~v3_1517448501_2599;
   assign v3_1517448501_2602 = f099 & v3_1517448501_2211;
   assign v3_1517448501_2603 = ~v3_1517448501_2604;
   assign v3_1517448501_2604 = ~v3_1517448501_2600 & ~v3_1517448501_2602;
   assign v3_1517448501_2605 = f100 & v3_1517448501_2213;
   assign v3_1517448501_2606 = ~v3_1517448501_2607;
   assign v3_1517448501_2607 = ~v3_1517448501_2603 & ~v3_1517448501_2605;
   assign v3_1517448501_2608 = f101 & v3_1517448501_2215;
   assign v3_1517448501_2609 = ~v3_1517448501_2610;
   assign v3_1517448501_2610 = ~v3_1517448501_2606 & ~v3_1517448501_2608;
   assign v3_1517448501_2611 = f102 & v3_1517448501_2217;
   assign v3_1517448501_2612 = ~v3_1517448501_2613;
   assign v3_1517448501_2613 = ~v3_1517448501_2609 & ~v3_1517448501_2611;
   assign v3_1517448501_2614 = f103 & v3_1517448501_2219;
   assign v3_1517448501_2615 = ~v3_1517448501_2616;
   assign v3_1517448501_2616 = ~v3_1517448501_2612 & ~v3_1517448501_2614;
   assign v3_1517448501_2617 = f104 & v3_1517448501_2221;
   assign v3_1517448501_2618 = ~v3_1517448501_2619;
   assign v3_1517448501_2619 = ~v3_1517448501_2615 & ~v3_1517448501_2617;
   assign v3_1517448501_2620 = f105 & v3_1517448501_2223;
   assign v3_1517448501_2621 = ~v3_1517448501_2622;
   assign v3_1517448501_2622 = ~v3_1517448501_2618 & ~v3_1517448501_2620;
   assign v3_1517448501_2623 = f106 & v3_1517448501_2225;
   assign v3_1517448501_2624 = ~v3_1517448501_2625;
   assign v3_1517448501_2625 = ~v3_1517448501_2621 & ~v3_1517448501_2623;
   assign v3_1517448501_2626 = f107 & v3_1517448501_2227;
   assign v3_1517448501_2627 = ~v3_1517448501_2628;
   assign v3_1517448501_2628 = ~v3_1517448501_2624 & ~v3_1517448501_2626;
   assign v3_1517448501_2629 = f108 & v3_1517448501_2229;
   assign v3_1517448501_2630 = ~v3_1517448501_2631;
   assign v3_1517448501_2631 = ~v3_1517448501_2627 & ~v3_1517448501_2629;
   assign v3_1517448501_2632 = f109 & v3_1517448501_2231;
   assign v3_1517448501_2633 = ~v3_1517448501_2634;
   assign v3_1517448501_2634 = ~v3_1517448501_2630 & ~v3_1517448501_2632;
   assign v3_1517448501_2635 = f110 & v3_1517448501_2233;
   assign v3_1517448501_2636 = ~v3_1517448501_2637;
   assign v3_1517448501_2637 = ~v3_1517448501_2633 & ~v3_1517448501_2635;
   assign v3_1517448501_2638 = f111 & v3_1517448501_2235;
   assign v3_1517448501_2639 = ~v3_1517448501_2640;
   assign v3_1517448501_2640 = ~v3_1517448501_2636 & ~v3_1517448501_2638;
   assign v3_1517448501_2641 = f112 & v3_1517448501_2237;
   assign v3_1517448501_2642 = ~v3_1517448501_2643;
   assign v3_1517448501_2643 = ~v3_1517448501_2639 & ~v3_1517448501_2641;
   assign v3_1517448501_2644 = f113 & v3_1517448501_2239;
   assign v3_1517448501_2645 = ~v3_1517448501_2646;
   assign v3_1517448501_2646 = ~v3_1517448501_2642 & ~v3_1517448501_2644;
   assign v3_1517448501_2647 = f114 & v3_1517448501_2241;
   assign v3_1517448501_2648 = ~v3_1517448501_2649;
   assign v3_1517448501_2649 = ~v3_1517448501_2645 & ~v3_1517448501_2647;
   assign v3_1517448501_2650 = f115 & v3_1517448501_2243;
   assign v3_1517448501_2651 = ~v3_1517448501_2652;
   assign v3_1517448501_2652 = ~v3_1517448501_2648 & ~v3_1517448501_2650;
   assign v3_1517448501_2653 = f116 & v3_1517448501_2245;
   assign v3_1517448501_2654 = ~v3_1517448501_2655;
   assign v3_1517448501_2655 = ~v3_1517448501_2651 & ~v3_1517448501_2653;
   assign v3_1517448501_2656 = f117 & v3_1517448501_2247;
   assign v3_1517448501_2657 = ~v3_1517448501_2658;
   assign v3_1517448501_2658 = ~v3_1517448501_2654 & ~v3_1517448501_2656;
   assign v3_1517448501_2659 = f118 & v3_1517448501_2249;
   assign v3_1517448501_2660 = ~v3_1517448501_2661;
   assign v3_1517448501_2661 = ~v3_1517448501_2657 & ~v3_1517448501_2659;
   assign v3_1517448501_2662 = f119 & v3_1517448501_2251;
   assign v3_1517448501_2663 = ~v3_1517448501_2664;
   assign v3_1517448501_2664 = ~v3_1517448501_2660 & ~v3_1517448501_2662;
   assign v3_1517448501_2665 = f120 & v3_1517448501_2253;
   assign v3_1517448501_2666 = ~v3_1517448501_2667;
   assign v3_1517448501_2667 = ~v3_1517448501_2663 & ~v3_1517448501_2665;
   assign v3_1517448501_2668 = f121 & v3_1517448501_2255;
   assign v3_1517448501_2669 = ~v3_1517448501_2670;
   assign v3_1517448501_2670 = ~v3_1517448501_2666 & ~v3_1517448501_2668;
   assign v3_1517448501_2671 = f122 & v3_1517448501_2257;
   assign v3_1517448501_2672 = ~v3_1517448501_2673;
   assign v3_1517448501_2673 = ~v3_1517448501_2669 & ~v3_1517448501_2671;
   assign v3_1517448501_2674 = f123 & v3_1517448501_2259;
   assign v3_1517448501_2675 = ~v3_1517448501_2676;
   assign v3_1517448501_2676 = ~v3_1517448501_2672 & ~v3_1517448501_2674;
   assign v3_1517448501_2677 = f124 & v3_1517448501_2261;
   assign v3_1517448501_2678 = ~v3_1517448501_2679;
   assign v3_1517448501_2679 = ~v3_1517448501_2675 & ~v3_1517448501_2677;
   assign v3_1517448501_2680 = f125 & v3_1517448501_2263;
   assign v3_1517448501_2681 = ~v3_1517448501_2682;
   assign v3_1517448501_2682 = ~v3_1517448501_2678 & ~v3_1517448501_2680;
   assign v3_1517448501_2683 = f126 & v3_1517448501_2265;
   assign v3_1517448501_2684 = ~v3_1517448501_2685;
   assign v3_1517448501_2685 = ~v3_1517448501_2681 & ~v3_1517448501_2683;
   assign v3_1517448501_2686 = f127 & v3_1517448501_2267;
   assign v3_1517448501_2687 = ~v3_1517448501_2688;
   assign v3_1517448501_2688 = ~v3_1517448501_2684 & ~v3_1517448501_2686;
   assign v3_1517448501_2689 = f128 & v3_1517448501_2269;
   assign v3_1517448501_2690 = ~v3_1517448501_2691;
   assign v3_1517448501_2691 = ~v3_1517448501_2687 & ~v3_1517448501_2689;
   assign v3_1517448501_2692 = f129 & v3_1517448501_2271;
   assign v3_1517448501_2693 = ~v3_1517448501_2694;
   assign v3_1517448501_2694 = ~v3_1517448501_2690 & ~v3_1517448501_2692;
   assign v3_1517448501_2695 = f130 & v3_1517448501_2273;
   assign v3_1517448501_2696 = ~v3_1517448501_2697;
   assign v3_1517448501_2697 = ~v3_1517448501_2693 & ~v3_1517448501_2695;
   assign v3_1517448501_2698 = f131 & v3_1517448501_2275;
   assign v3_1517448501_2699 = ~v3_1517448501_2700;
   assign v3_1517448501_2700 = ~v3_1517448501_2696 & ~v3_1517448501_2698;
   assign v3_1517448501_2701 = f132 & v3_1517448501_2277;
   assign v3_1517448501_2702 = ~v3_1517448501_2703;
   assign v3_1517448501_2703 = ~v3_1517448501_2699 & ~v3_1517448501_2701;
   assign v3_1517448501_2704 = f133 & v3_1517448501_2279;
   assign v3_1517448501_2705 = ~v3_1517448501_2706;
   assign v3_1517448501_2706 = ~v3_1517448501_2702 & ~v3_1517448501_2704;
   assign v3_1517448501_2707 = f134 & v3_1517448501_2281;
   assign v3_1517448501_2708 = ~v3_1517448501_2709;
   assign v3_1517448501_2709 = ~v3_1517448501_2705 & ~v3_1517448501_2707;
   assign v3_1517448501_2710 = f135 & v3_1517448501_2283;
   assign v3_1517448501_2711 = ~v3_1517448501_2712;
   assign v3_1517448501_2712 = ~v3_1517448501_2708 & ~v3_1517448501_2710;
   assign v3_1517448501_2713 = f136 & v3_1517448501_2285;
   assign v3_1517448501_2714 = ~v3_1517448501_2715;
   assign v3_1517448501_2715 = ~v3_1517448501_2711 & ~v3_1517448501_2713;
   assign v3_1517448501_2716 = f137 & v3_1517448501_2287;
   assign v3_1517448501_2717 = ~v3_1517448501_2718;
   assign v3_1517448501_2718 = ~v3_1517448501_2714 & ~v3_1517448501_2716;
   assign v3_1517448501_2719 = f138 & v3_1517448501_2289;
   assign v3_1517448501_2720 = ~v3_1517448501_2721;
   assign v3_1517448501_2721 = ~v3_1517448501_2717 & ~v3_1517448501_2719;
   assign v3_1517448501_2722 = f139 & v3_1517448501_2291;
   assign v3_1517448501_2723 = ~v3_1517448501_2724;
   assign v3_1517448501_2724 = ~v3_1517448501_2720 & ~v3_1517448501_2722;
   assign v3_1517448501_2725 = f140 & v3_1517448501_2293;
   assign v3_1517448501_2726 = ~v3_1517448501_2727;
   assign v3_1517448501_2727 = ~v3_1517448501_2723 & ~v3_1517448501_2725;
   assign v3_1517448501_2728 = f141 & v3_1517448501_2295;
   assign v3_1517448501_2729 = ~v3_1517448501_2730;
   assign v3_1517448501_2730 = ~v3_1517448501_2726 & ~v3_1517448501_2728;
   assign v3_1517448501_2731 = f142 & v3_1517448501_2297;
   assign v3_1517448501_2732 = ~v3_1517448501_2733;
   assign v3_1517448501_2733 = ~v3_1517448501_2729 & ~v3_1517448501_2731;
   assign v3_1517448501_2734 = f143 & v3_1517448501_2299;
   assign v3_1517448501_2735 = ~v3_1517448501_2736;
   assign v3_1517448501_2736 = ~v3_1517448501_2732 & ~v3_1517448501_2734;
   assign v3_1517448501_2737 = f144 & v3_1517448501_2301;
   assign v3_1517448501_2738 = ~v3_1517448501_2739;
   assign v3_1517448501_2739 = ~v3_1517448501_2735 & ~v3_1517448501_2737;
   assign v3_1517448501_2740 = f145 & v3_1517448501_2303;
   assign v3_1517448501_2741 = ~v3_1517448501_2742;
   assign v3_1517448501_2742 = ~v3_1517448501_2738 & ~v3_1517448501_2740;
   assign v3_1517448501_2743 = f146 & v3_1517448501_2305;
   assign v3_1517448501_2744 = ~v3_1517448501_2745;
   assign v3_1517448501_2745 = ~v3_1517448501_2741 & ~v3_1517448501_2743;
   assign v3_1517448501_2746 = v3_1517448501_2309 & ~v3_1517448501_2744;
   assign v3_1517448501_2747 = ~a_start_initiator_0 & a_wait_resp_initiator_0;
   assign v3_1517448501_2748 = ~v3_1517448501_2749;
   assign v3_1517448501_2749 = a_start_initiator_0 & ~a_wait_resp_initiator_0;
   assign v3_1517448501_2750 = a_got_resp_initiator_0 & v3_1517448501_2748;
   assign v3_1517448501_2751 = ~v3_1517448501_2752;
   assign v3_1517448501_2752 = ~v3_1517448501_2747 & ~v3_1517448501_2750;
   assign v3_1517448501_2753 = ~v3_1517448501_2754;
   assign v3_1517448501_2754 = ~a_got_resp_initiator_0 & ~v3_1517448501_2748;
   assign v3_1517448501_2755 = a_commited_initiator_0 & v3_1517448501_2753;
   assign v3_1517448501_2756 = ~v3_1517448501_2757;
   assign v3_1517448501_2757 = ~v3_1517448501_2751 & ~v3_1517448501_2755;
   assign v3_1517448501_2758 = ~v3_1517448501_2759;
   assign v3_1517448501_2759 = ~a_commited_initiator_0 & ~v3_1517448501_2753;
   assign v3_1517448501_2760 = a_finished_initiator_0 & v3_1517448501_2758;
   assign v3_1517448501_2761 = ~v3_1517448501_2762;
   assign v3_1517448501_2762 = ~v3_1517448501_2756 & ~v3_1517448501_2760;
   assign v3_1517448501_2763 = ~v3_1517448501_2764;
   assign v3_1517448501_2764 = ~a_finished_initiator_0 & ~v3_1517448501_2758;
   assign v3_1517448501_2765 = a_corrupted_initiator_0 & v3_1517448501_2763;
   assign v3_1517448501_2766 = ~v3_1517448501_2767;
   assign v3_1517448501_2767 = ~v3_1517448501_2761 & ~v3_1517448501_2765;
   assign v3_1517448501_2768 = ~v3_1517448501_2769;
   assign v3_1517448501_2769 = ~a_corrupted_initiator_0 & ~v3_1517448501_2763;
   assign v3_1517448501_2770 = ~v3_1517448501_2766 & v3_1517448501_2768;
   assign v3_1517448501_2771 = ~a_start_initiator_1 & a_wait_resp_initiator_1;
   assign v3_1517448501_2772 = ~v3_1517448501_2773;
   assign v3_1517448501_2773 = a_start_initiator_1 & ~a_wait_resp_initiator_1;
   assign v3_1517448501_2774 = a_got_resp_initiator_1 & v3_1517448501_2772;
   assign v3_1517448501_2775 = ~v3_1517448501_2776;
   assign v3_1517448501_2776 = ~v3_1517448501_2771 & ~v3_1517448501_2774;
   assign v3_1517448501_2777 = ~v3_1517448501_2778;
   assign v3_1517448501_2778 = ~a_got_resp_initiator_1 & ~v3_1517448501_2772;
   assign v3_1517448501_2779 = a_commited_initiator_1 & v3_1517448501_2777;
   assign v3_1517448501_2780 = ~v3_1517448501_2781;
   assign v3_1517448501_2781 = ~v3_1517448501_2775 & ~v3_1517448501_2779;
   assign v3_1517448501_2782 = ~v3_1517448501_2783;
   assign v3_1517448501_2783 = ~a_commited_initiator_1 & ~v3_1517448501_2777;
   assign v3_1517448501_2784 = a_finished_initiator_1 & v3_1517448501_2782;
   assign v3_1517448501_2785 = ~v3_1517448501_2786;
   assign v3_1517448501_2786 = ~v3_1517448501_2780 & ~v3_1517448501_2784;
   assign v3_1517448501_2787 = ~v3_1517448501_2788;
   assign v3_1517448501_2788 = ~a_finished_initiator_1 & ~v3_1517448501_2782;
   assign v3_1517448501_2789 = a_corrupted_initiator_1 & v3_1517448501_2787;
   assign v3_1517448501_2790 = ~v3_1517448501_2791;
   assign v3_1517448501_2791 = ~v3_1517448501_2785 & ~v3_1517448501_2789;
   assign v3_1517448501_2792 = v3_1517448501_2770 & ~v3_1517448501_2790;
   assign v3_1517448501_2793 = ~v3_1517448501_2794;
   assign v3_1517448501_2794 = ~a_corrupted_initiator_1 & ~v3_1517448501_2787;
   assign v3_1517448501_2795 = v3_1517448501_2792 & v3_1517448501_2793;
   assign v3_1517448501_2796 = ~a_start_initiator_2 & a_wait_resp_initiator_2;
   assign v3_1517448501_2797 = ~v3_1517448501_2798;
   assign v3_1517448501_2798 = a_start_initiator_2 & ~a_wait_resp_initiator_2;
   assign v3_1517448501_2799 = a_got_resp_initiator_2 & v3_1517448501_2797;
   assign v3_1517448501_2800 = ~v3_1517448501_2801;
   assign v3_1517448501_2801 = ~v3_1517448501_2796 & ~v3_1517448501_2799;
   assign v3_1517448501_2802 = ~v3_1517448501_2803;
   assign v3_1517448501_2803 = ~a_got_resp_initiator_2 & ~v3_1517448501_2797;
   assign v3_1517448501_2804 = a_commited_initiator_2 & v3_1517448501_2802;
   assign v3_1517448501_2805 = ~v3_1517448501_2806;
   assign v3_1517448501_2806 = ~v3_1517448501_2800 & ~v3_1517448501_2804;
   assign v3_1517448501_2807 = ~v3_1517448501_2808;
   assign v3_1517448501_2808 = ~a_commited_initiator_2 & ~v3_1517448501_2802;
   assign v3_1517448501_2809 = a_finished_initiator_2 & v3_1517448501_2807;
   assign v3_1517448501_2810 = ~v3_1517448501_2811;
   assign v3_1517448501_2811 = ~v3_1517448501_2805 & ~v3_1517448501_2809;
   assign v3_1517448501_2812 = ~v3_1517448501_2813;
   assign v3_1517448501_2813 = ~a_finished_initiator_2 & ~v3_1517448501_2807;
   assign v3_1517448501_2814 = a_corrupted_initiator_2 & v3_1517448501_2812;
   assign v3_1517448501_2815 = ~v3_1517448501_2816;
   assign v3_1517448501_2816 = ~v3_1517448501_2810 & ~v3_1517448501_2814;
   assign v3_1517448501_2817 = v3_1517448501_2795 & ~v3_1517448501_2815;
   assign v3_1517448501_2818 = ~v3_1517448501_2819;
   assign v3_1517448501_2819 = ~a_corrupted_initiator_2 & ~v3_1517448501_2812;
   assign v3_1517448501_2820 = v3_1517448501_2817 & v3_1517448501_2818;
   assign v3_1517448501_2821 = ~a_start_responder_0 & a_got_msg_responder_0;
   assign v3_1517448501_2822 = ~v3_1517448501_2823;
   assign v3_1517448501_2823 = a_start_responder_0 & ~a_got_msg_responder_0;
   assign v3_1517448501_2824 = a_send_reply_responder_0 & v3_1517448501_2822;
   assign v3_1517448501_2825 = ~v3_1517448501_2826;
   assign v3_1517448501_2826 = ~v3_1517448501_2821 & ~v3_1517448501_2824;
   assign v3_1517448501_2827 = ~v3_1517448501_2828;
   assign v3_1517448501_2828 = ~a_send_reply_responder_0 & ~v3_1517448501_2822;
   assign v3_1517448501_2829 = a_wait_resp_responder_0 & v3_1517448501_2827;
   assign v3_1517448501_2830 = ~v3_1517448501_2831;
   assign v3_1517448501_2831 = ~v3_1517448501_2825 & ~v3_1517448501_2829;
   assign v3_1517448501_2832 = ~v3_1517448501_2833;
   assign v3_1517448501_2833 = ~a_wait_resp_responder_0 & ~v3_1517448501_2827;
   assign v3_1517448501_2834 = a_got_resp_responder_0 & v3_1517448501_2832;
   assign v3_1517448501_2835 = ~v3_1517448501_2836;
   assign v3_1517448501_2836 = ~v3_1517448501_2830 & ~v3_1517448501_2834;
   assign v3_1517448501_2837 = ~v3_1517448501_2838;
   assign v3_1517448501_2838 = ~a_got_resp_responder_0 & ~v3_1517448501_2832;
   assign v3_1517448501_2839 = a_finished_responder_0 & v3_1517448501_2837;
   assign v3_1517448501_2840 = ~v3_1517448501_2841;
   assign v3_1517448501_2841 = ~v3_1517448501_2835 & ~v3_1517448501_2839;
   assign v3_1517448501_2842 = ~v3_1517448501_2843;
   assign v3_1517448501_2843 = ~a_finished_responder_0 & ~v3_1517448501_2837;
   assign v3_1517448501_2844 = a_corrupted_responder_0 & v3_1517448501_2842;
   assign v3_1517448501_2845 = ~v3_1517448501_2846;
   assign v3_1517448501_2846 = ~v3_1517448501_2840 & ~v3_1517448501_2844;
   assign v3_1517448501_2847 = v3_1517448501_2820 & ~v3_1517448501_2845;
   assign v3_1517448501_2848 = ~v3_1517448501_2849;
   assign v3_1517448501_2849 = ~a_corrupted_responder_0 & ~v3_1517448501_2842;
   assign v3_1517448501_2850 = v3_1517448501_2847 & v3_1517448501_2848;
   assign v3_1517448501_2851 = ~a_start_responder_1 & a_got_msg_responder_1;
   assign v3_1517448501_2852 = ~v3_1517448501_2853;
   assign v3_1517448501_2853 = a_start_responder_1 & ~a_got_msg_responder_1;
   assign v3_1517448501_2854 = a_send_reply_responder_1 & v3_1517448501_2852;
   assign v3_1517448501_2855 = ~v3_1517448501_2856;
   assign v3_1517448501_2856 = ~v3_1517448501_2851 & ~v3_1517448501_2854;
   assign v3_1517448501_2857 = ~v3_1517448501_2858;
   assign v3_1517448501_2858 = ~a_send_reply_responder_1 & ~v3_1517448501_2852;
   assign v3_1517448501_2859 = a_wait_resp_responder_1 & v3_1517448501_2857;
   assign v3_1517448501_2860 = ~v3_1517448501_2861;
   assign v3_1517448501_2861 = ~v3_1517448501_2855 & ~v3_1517448501_2859;
   assign v3_1517448501_2862 = ~v3_1517448501_2863;
   assign v3_1517448501_2863 = ~a_wait_resp_responder_1 & ~v3_1517448501_2857;
   assign v3_1517448501_2864 = a_got_resp_responder_1 & v3_1517448501_2862;
   assign v3_1517448501_2865 = ~v3_1517448501_2866;
   assign v3_1517448501_2866 = ~v3_1517448501_2860 & ~v3_1517448501_2864;
   assign v3_1517448501_2867 = ~v3_1517448501_2868;
   assign v3_1517448501_2868 = ~a_got_resp_responder_1 & ~v3_1517448501_2862;
   assign v3_1517448501_2869 = a_finished_responder_1 & v3_1517448501_2867;
   assign v3_1517448501_2870 = ~v3_1517448501_2871;
   assign v3_1517448501_2871 = ~v3_1517448501_2865 & ~v3_1517448501_2869;
   assign v3_1517448501_2872 = ~v3_1517448501_2873;
   assign v3_1517448501_2873 = ~a_finished_responder_1 & ~v3_1517448501_2867;
   assign v3_1517448501_2874 = a_corrupted_responder_1 & v3_1517448501_2872;
   assign v3_1517448501_2875 = ~v3_1517448501_2876;
   assign v3_1517448501_2876 = ~v3_1517448501_2870 & ~v3_1517448501_2874;
   assign v3_1517448501_2877 = v3_1517448501_2850 & ~v3_1517448501_2875;
   assign v3_1517448501_2878 = ~v3_1517448501_2879;
   assign v3_1517448501_2879 = ~a_corrupted_responder_1 & ~v3_1517448501_2872;
   assign v3_1517448501_2880 = v3_1517448501_2877 & v3_1517448501_2878;
   assign v3_1517448501_2881 = ~a_start_responder_2 & a_got_msg_responder_2;
   assign v3_1517448501_2882 = ~v3_1517448501_2883;
   assign v3_1517448501_2883 = a_start_responder_2 & ~a_got_msg_responder_2;
   assign v3_1517448501_2884 = a_send_reply_responder_2 & v3_1517448501_2882;
   assign v3_1517448501_2885 = ~v3_1517448501_2886;
   assign v3_1517448501_2886 = ~v3_1517448501_2881 & ~v3_1517448501_2884;
   assign v3_1517448501_2887 = ~v3_1517448501_2888;
   assign v3_1517448501_2888 = ~a_send_reply_responder_2 & ~v3_1517448501_2882;
   assign v3_1517448501_2889 = a_wait_resp_responder_2 & v3_1517448501_2887;
   assign v3_1517448501_2890 = ~v3_1517448501_2891;
   assign v3_1517448501_2891 = ~v3_1517448501_2885 & ~v3_1517448501_2889;
   assign v3_1517448501_2892 = ~v3_1517448501_2893;
   assign v3_1517448501_2893 = ~a_wait_resp_responder_2 & ~v3_1517448501_2887;
   assign v3_1517448501_2894 = a_got_resp_responder_2 & v3_1517448501_2892;
   assign v3_1517448501_2895 = ~v3_1517448501_2896;
   assign v3_1517448501_2896 = ~v3_1517448501_2890 & ~v3_1517448501_2894;
   assign v3_1517448501_2897 = ~v3_1517448501_2898;
   assign v3_1517448501_2898 = ~a_got_resp_responder_2 & ~v3_1517448501_2892;
   assign v3_1517448501_2899 = a_finished_responder_2 & v3_1517448501_2897;
   assign v3_1517448501_2900 = ~v3_1517448501_2901;
   assign v3_1517448501_2901 = ~v3_1517448501_2895 & ~v3_1517448501_2899;
   assign v3_1517448501_2902 = ~v3_1517448501_2903;
   assign v3_1517448501_2903 = ~a_finished_responder_2 & ~v3_1517448501_2897;
   assign v3_1517448501_2904 = a_corrupted_responder_2 & v3_1517448501_2902;
   assign v3_1517448501_2905 = ~v3_1517448501_2906;
   assign v3_1517448501_2906 = ~v3_1517448501_2900 & ~v3_1517448501_2904;
   assign v3_1517448501_2907 = v3_1517448501_2880 & ~v3_1517448501_2905;
   assign v3_1517448501_2908 = ~v3_1517448501_2909;
   assign v3_1517448501_2909 = ~a_corrupted_responder_2 & ~v3_1517448501_2902;
   assign v3_1517448501_2910 = v3_1517448501_2907 & v3_1517448501_2908;
   assign v3_1517448501_2911 = ~a_q & a_got3;
   assign v3_1517448501_2912 = ~v3_1517448501_2913;
   assign v3_1517448501_2913 = a_q & ~a_got3;
   assign v3_1517448501_2914 = a_c1 & v3_1517448501_2912;
   assign v3_1517448501_2915 = ~v3_1517448501_2916;
   assign v3_1517448501_2916 = ~v3_1517448501_2911 & ~v3_1517448501_2914;
   assign v3_1517448501_2917 = ~v3_1517448501_2918;
   assign v3_1517448501_2918 = ~a_c1 & ~v3_1517448501_2912;
   assign v3_1517448501_2919 = a_c2 & v3_1517448501_2917;
   assign v3_1517448501_2920 = ~v3_1517448501_2921;
   assign v3_1517448501_2921 = ~v3_1517448501_2915 & ~v3_1517448501_2919;
   assign v3_1517448501_2922 = ~v3_1517448501_2923;
   assign v3_1517448501_2923 = ~a_c2 & ~v3_1517448501_2917;
   assign v3_1517448501_2924 = a_d1 & v3_1517448501_2922;
   assign v3_1517448501_2925 = ~v3_1517448501_2926;
   assign v3_1517448501_2926 = ~v3_1517448501_2920 & ~v3_1517448501_2924;
   assign v3_1517448501_2927 = ~v3_1517448501_2928;
   assign v3_1517448501_2928 = ~a_d1 & ~v3_1517448501_2922;
   assign v3_1517448501_2929 = a_got2 & v3_1517448501_2927;
   assign v3_1517448501_2930 = ~v3_1517448501_2931;
   assign v3_1517448501_2931 = ~v3_1517448501_2925 & ~v3_1517448501_2929;
   assign v3_1517448501_2932 = ~v3_1517448501_2933;
   assign v3_1517448501_2933 = ~a_got2 & ~v3_1517448501_2927;
   assign v3_1517448501_2934 = a_e1 & v3_1517448501_2932;
   assign v3_1517448501_2935 = ~v3_1517448501_2936;
   assign v3_1517448501_2936 = ~v3_1517448501_2930 & ~v3_1517448501_2934;
   assign v3_1517448501_2937 = ~v3_1517448501_2938;
   assign v3_1517448501_2938 = ~a_e1 & ~v3_1517448501_2932;
   assign v3_1517448501_2939 = a_f1 & v3_1517448501_2937;
   assign v3_1517448501_2940 = ~v3_1517448501_2941;
   assign v3_1517448501_2941 = ~v3_1517448501_2935 & ~v3_1517448501_2939;
   assign v3_1517448501_2942 = v3_1517448501_2910 & ~v3_1517448501_2940;
   assign v3_1517448501_2943 = ~v3_1517448501_2944;
   assign v3_1517448501_2944 = ~a_f1 & ~v3_1517448501_2937;
   assign v3_1517448501_2945 = v3_1517448501_2942 & v3_1517448501_2943;
   assign v3_1517448501_2946 = v3_1517448501_2746 & v3_1517448501_2945;
   assign v3_1517448501_2947 = v3_1517448501_650 & v3_1517448501_665;
   assign v3_1517448501_2948 = ~v3_1517448501_2949;
   assign v3_1517448501_2949 = ~v3_1517448501_650 & ~v3_1517448501_665;
   assign v3_1517448501_2950 = v3_1517448501_680 & v3_1517448501_2948;
   assign v3_1517448501_2951 = ~v3_1517448501_2952;
   assign v3_1517448501_2952 = ~v3_1517448501_2947 & ~v3_1517448501_2950;
   assign v3_1517448501_2953 = ~v3_1517448501_2954;
   assign v3_1517448501_2954 = ~v3_1517448501_680 & ~v3_1517448501_2948;
   assign v3_1517448501_2955 = v3_1517448501_688 & v3_1517448501_2953;
   assign v3_1517448501_2956 = ~v3_1517448501_2957;
   assign v3_1517448501_2957 = ~v3_1517448501_2951 & ~v3_1517448501_2955;
   assign v3_1517448501_2958 = ~v3_1517448501_2959;
   assign v3_1517448501_2959 = ~v3_1517448501_688 & ~v3_1517448501_2953;
   assign v3_1517448501_2960 = v3_1517448501_696 & v3_1517448501_2958;
   assign v3_1517448501_2961 = ~v3_1517448501_2962;
   assign v3_1517448501_2962 = ~v3_1517448501_2956 & ~v3_1517448501_2960;
   assign v3_1517448501_2963 = ~v3_1517448501_2964;
   assign v3_1517448501_2964 = ~v3_1517448501_696 & ~v3_1517448501_2958;
   assign v3_1517448501_2965 = v3_1517448501_699 & v3_1517448501_2963;
   assign v3_1517448501_2966 = ~v3_1517448501_2967;
   assign v3_1517448501_2967 = ~v3_1517448501_2961 & ~v3_1517448501_2965;
   assign v3_1517448501_2968 = ~v3_1517448501_2969;
   assign v3_1517448501_2969 = ~v3_1517448501_699 & ~v3_1517448501_2963;
   assign v3_1517448501_2970 = ~v3_1517448501_2966 & v3_1517448501_2968;
   assign v3_1517448501_2971 = v3_1517448501_705 & v3_1517448501_720;
   assign v3_1517448501_2972 = ~v3_1517448501_2973;
   assign v3_1517448501_2973 = ~v3_1517448501_705 & ~v3_1517448501_720;
   assign v3_1517448501_2974 = v3_1517448501_735 & v3_1517448501_2972;
   assign v3_1517448501_2975 = ~v3_1517448501_2976;
   assign v3_1517448501_2976 = ~v3_1517448501_2971 & ~v3_1517448501_2974;
   assign v3_1517448501_2977 = ~v3_1517448501_2978;
   assign v3_1517448501_2978 = ~v3_1517448501_735 & ~v3_1517448501_2972;
   assign v3_1517448501_2979 = v3_1517448501_743 & v3_1517448501_2977;
   assign v3_1517448501_2980 = ~v3_1517448501_2981;
   assign v3_1517448501_2981 = ~v3_1517448501_2975 & ~v3_1517448501_2979;
   assign v3_1517448501_2982 = ~v3_1517448501_2983;
   assign v3_1517448501_2983 = ~v3_1517448501_743 & ~v3_1517448501_2977;
   assign v3_1517448501_2984 = v3_1517448501_751 & v3_1517448501_2982;
   assign v3_1517448501_2985 = ~v3_1517448501_2986;
   assign v3_1517448501_2986 = ~v3_1517448501_2980 & ~v3_1517448501_2984;
   assign v3_1517448501_2987 = ~v3_1517448501_2988;
   assign v3_1517448501_2988 = ~v3_1517448501_751 & ~v3_1517448501_2982;
   assign v3_1517448501_2989 = v3_1517448501_754 & v3_1517448501_2987;
   assign v3_1517448501_2990 = ~v3_1517448501_2991;
   assign v3_1517448501_2991 = ~v3_1517448501_2985 & ~v3_1517448501_2989;
   assign v3_1517448501_2992 = v3_1517448501_2970 & ~v3_1517448501_2990;
   assign v3_1517448501_2993 = ~v3_1517448501_2994;
   assign v3_1517448501_2994 = ~v3_1517448501_754 & ~v3_1517448501_2987;
   assign v3_1517448501_2995 = v3_1517448501_2992 & v3_1517448501_2993;
   assign v3_1517448501_2996 = v3_1517448501_760 & v3_1517448501_775;
   assign v3_1517448501_2997 = ~v3_1517448501_2998;
   assign v3_1517448501_2998 = ~v3_1517448501_760 & ~v3_1517448501_775;
   assign v3_1517448501_2999 = v3_1517448501_790 & v3_1517448501_2997;
   assign v3_1517448501_3000 = ~v3_1517448501_3001;
   assign v3_1517448501_3001 = ~v3_1517448501_2996 & ~v3_1517448501_2999;
   assign v3_1517448501_3002 = ~v3_1517448501_3003;
   assign v3_1517448501_3003 = ~v3_1517448501_790 & ~v3_1517448501_2997;
   assign v3_1517448501_3004 = v3_1517448501_798 & v3_1517448501_3002;
   assign v3_1517448501_3005 = ~v3_1517448501_3006;
   assign v3_1517448501_3006 = ~v3_1517448501_3000 & ~v3_1517448501_3004;
   assign v3_1517448501_3007 = ~v3_1517448501_3008;
   assign v3_1517448501_3008 = ~v3_1517448501_798 & ~v3_1517448501_3002;
   assign v3_1517448501_3009 = v3_1517448501_806 & v3_1517448501_3007;
   assign v3_1517448501_3010 = ~v3_1517448501_3011;
   assign v3_1517448501_3011 = ~v3_1517448501_3005 & ~v3_1517448501_3009;
   assign v3_1517448501_3012 = ~v3_1517448501_3013;
   assign v3_1517448501_3013 = ~v3_1517448501_806 & ~v3_1517448501_3007;
   assign v3_1517448501_3014 = v3_1517448501_809 & v3_1517448501_3012;
   assign v3_1517448501_3015 = ~v3_1517448501_3016;
   assign v3_1517448501_3016 = ~v3_1517448501_3010 & ~v3_1517448501_3014;
   assign v3_1517448501_3017 = v3_1517448501_2995 & ~v3_1517448501_3015;
   assign v3_1517448501_3018 = ~v3_1517448501_3019;
   assign v3_1517448501_3019 = ~v3_1517448501_809 & ~v3_1517448501_3012;
   assign v3_1517448501_3020 = v3_1517448501_3017 & v3_1517448501_3018;
   assign v3_1517448501_3021 = v3_1517448501_835 & v3_1517448501_886;
   assign v3_1517448501_3022 = ~v3_1517448501_3023;
   assign v3_1517448501_3023 = ~v3_1517448501_835 & ~v3_1517448501_886;
   assign v3_1517448501_3024 = v3_1517448501_894 & v3_1517448501_3022;
   assign v3_1517448501_3025 = ~v3_1517448501_3026;
   assign v3_1517448501_3026 = ~v3_1517448501_3021 & ~v3_1517448501_3024;
   assign v3_1517448501_3027 = ~v3_1517448501_3028;
   assign v3_1517448501_3028 = ~v3_1517448501_894 & ~v3_1517448501_3022;
   assign v3_1517448501_3029 = v3_1517448501_907 & v3_1517448501_3027;
   assign v3_1517448501_3030 = ~v3_1517448501_3031;
   assign v3_1517448501_3031 = ~v3_1517448501_3025 & ~v3_1517448501_3029;
   assign v3_1517448501_3032 = ~v3_1517448501_3033;
   assign v3_1517448501_3033 = ~v3_1517448501_907 & ~v3_1517448501_3027;
   assign v3_1517448501_3034 = v3_1517448501_919 & v3_1517448501_3032;
   assign v3_1517448501_3035 = ~v3_1517448501_3036;
   assign v3_1517448501_3036 = ~v3_1517448501_3030 & ~v3_1517448501_3034;
   assign v3_1517448501_3037 = ~v3_1517448501_3038;
   assign v3_1517448501_3038 = ~v3_1517448501_919 & ~v3_1517448501_3032;
   assign v3_1517448501_3039 = v3_1517448501_922 & v3_1517448501_3037;
   assign v3_1517448501_3040 = ~v3_1517448501_3041;
   assign v3_1517448501_3041 = ~v3_1517448501_3035 & ~v3_1517448501_3039;
   assign v3_1517448501_3042 = ~v3_1517448501_3043;
   assign v3_1517448501_3043 = ~v3_1517448501_922 & ~v3_1517448501_3037;
   assign v3_1517448501_3044 = v3_1517448501_927 & v3_1517448501_3042;
   assign v3_1517448501_3045 = ~v3_1517448501_3046;
   assign v3_1517448501_3046 = ~v3_1517448501_3040 & ~v3_1517448501_3044;
   assign v3_1517448501_3047 = v3_1517448501_3020 & ~v3_1517448501_3045;
   assign v3_1517448501_3048 = ~v3_1517448501_3049;
   assign v3_1517448501_3049 = ~v3_1517448501_927 & ~v3_1517448501_3042;
   assign v3_1517448501_3050 = v3_1517448501_3047 & v3_1517448501_3048;
   assign v3_1517448501_3051 = v3_1517448501_953 & v3_1517448501_1004;
   assign v3_1517448501_3052 = ~v3_1517448501_3053;
   assign v3_1517448501_3053 = ~v3_1517448501_953 & ~v3_1517448501_1004;
   assign v3_1517448501_3054 = v3_1517448501_1012 & v3_1517448501_3052;
   assign v3_1517448501_3055 = ~v3_1517448501_3056;
   assign v3_1517448501_3056 = ~v3_1517448501_3051 & ~v3_1517448501_3054;
   assign v3_1517448501_3057 = ~v3_1517448501_3058;
   assign v3_1517448501_3058 = ~v3_1517448501_1012 & ~v3_1517448501_3052;
   assign v3_1517448501_3059 = v3_1517448501_1025 & v3_1517448501_3057;
   assign v3_1517448501_3060 = ~v3_1517448501_3061;
   assign v3_1517448501_3061 = ~v3_1517448501_3055 & ~v3_1517448501_3059;
   assign v3_1517448501_3062 = ~v3_1517448501_3063;
   assign v3_1517448501_3063 = ~v3_1517448501_1025 & ~v3_1517448501_3057;
   assign v3_1517448501_3064 = v3_1517448501_1037 & v3_1517448501_3062;
   assign v3_1517448501_3065 = ~v3_1517448501_3066;
   assign v3_1517448501_3066 = ~v3_1517448501_3060 & ~v3_1517448501_3064;
   assign v3_1517448501_3067 = ~v3_1517448501_3068;
   assign v3_1517448501_3068 = ~v3_1517448501_1037 & ~v3_1517448501_3062;
   assign v3_1517448501_3069 = v3_1517448501_1040 & v3_1517448501_3067;
   assign v3_1517448501_3070 = ~v3_1517448501_3071;
   assign v3_1517448501_3071 = ~v3_1517448501_3065 & ~v3_1517448501_3069;
   assign v3_1517448501_3072 = ~v3_1517448501_3073;
   assign v3_1517448501_3073 = ~v3_1517448501_1040 & ~v3_1517448501_3067;
   assign v3_1517448501_3074 = v3_1517448501_1045 & v3_1517448501_3072;
   assign v3_1517448501_3075 = ~v3_1517448501_3076;
   assign v3_1517448501_3076 = ~v3_1517448501_3070 & ~v3_1517448501_3074;
   assign v3_1517448501_3077 = v3_1517448501_3050 & ~v3_1517448501_3075;
   assign v3_1517448501_3078 = ~v3_1517448501_3079;
   assign v3_1517448501_3079 = ~v3_1517448501_1045 & ~v3_1517448501_3072;
   assign v3_1517448501_3080 = v3_1517448501_3077 & v3_1517448501_3078;
   assign v3_1517448501_3081 = v3_1517448501_1071 & v3_1517448501_1122;
   assign v3_1517448501_3082 = ~v3_1517448501_3083;
   assign v3_1517448501_3083 = ~v3_1517448501_1071 & ~v3_1517448501_1122;
   assign v3_1517448501_3084 = v3_1517448501_1130 & v3_1517448501_3082;
   assign v3_1517448501_3085 = ~v3_1517448501_3086;
   assign v3_1517448501_3086 = ~v3_1517448501_3081 & ~v3_1517448501_3084;
   assign v3_1517448501_3087 = ~v3_1517448501_3088;
   assign v3_1517448501_3088 = ~v3_1517448501_1130 & ~v3_1517448501_3082;
   assign v3_1517448501_3089 = v3_1517448501_1143 & v3_1517448501_3087;
   assign v3_1517448501_3090 = ~v3_1517448501_3091;
   assign v3_1517448501_3091 = ~v3_1517448501_3085 & ~v3_1517448501_3089;
   assign v3_1517448501_3092 = ~v3_1517448501_3093;
   assign v3_1517448501_3093 = ~v3_1517448501_1143 & ~v3_1517448501_3087;
   assign v3_1517448501_3094 = v3_1517448501_1155 & v3_1517448501_3092;
   assign v3_1517448501_3095 = ~v3_1517448501_3096;
   assign v3_1517448501_3096 = ~v3_1517448501_3090 & ~v3_1517448501_3094;
   assign v3_1517448501_3097 = ~v3_1517448501_3098;
   assign v3_1517448501_3098 = ~v3_1517448501_1155 & ~v3_1517448501_3092;
   assign v3_1517448501_3099 = v3_1517448501_1158 & v3_1517448501_3097;
   assign v3_1517448501_3100 = ~v3_1517448501_3101;
   assign v3_1517448501_3101 = ~v3_1517448501_3095 & ~v3_1517448501_3099;
   assign v3_1517448501_3102 = ~v3_1517448501_3103;
   assign v3_1517448501_3103 = ~v3_1517448501_1158 & ~v3_1517448501_3097;
   assign v3_1517448501_3104 = v3_1517448501_1163 & v3_1517448501_3102;
   assign v3_1517448501_3105 = ~v3_1517448501_3106;
   assign v3_1517448501_3106 = ~v3_1517448501_3100 & ~v3_1517448501_3104;
   assign v3_1517448501_3107 = v3_1517448501_3080 & ~v3_1517448501_3105;
   assign v3_1517448501_3108 = ~v3_1517448501_3109;
   assign v3_1517448501_3109 = ~v3_1517448501_1163 & ~v3_1517448501_3102;
   assign v3_1517448501_3110 = v3_1517448501_3107 & v3_1517448501_3108;
   assign v3_1517448501_3111 = v3_1517448501_1218 & v3_1517448501_1201;
   assign v3_1517448501_3112 = ~v3_1517448501_3113;
   assign v3_1517448501_3113 = ~v3_1517448501_1218 & ~v3_1517448501_1201;
   assign v3_1517448501_3114 = v3_1517448501_1226 & v3_1517448501_3112;
   assign v3_1517448501_3115 = ~v3_1517448501_3116;
   assign v3_1517448501_3116 = ~v3_1517448501_3111 & ~v3_1517448501_3114;
   assign v3_1517448501_3117 = ~v3_1517448501_3118;
   assign v3_1517448501_3118 = ~v3_1517448501_1226 & ~v3_1517448501_3112;
   assign v3_1517448501_3119 = v3_1517448501_1235 & v3_1517448501_3117;
   assign v3_1517448501_3120 = ~v3_1517448501_3121;
   assign v3_1517448501_3121 = ~v3_1517448501_3115 & ~v3_1517448501_3119;
   assign v3_1517448501_3122 = ~v3_1517448501_3123;
   assign v3_1517448501_3123 = ~v3_1517448501_1235 & ~v3_1517448501_3117;
   assign v3_1517448501_3124 = v3_1517448501_1241 & v3_1517448501_3122;
   assign v3_1517448501_3125 = ~v3_1517448501_3126;
   assign v3_1517448501_3126 = ~v3_1517448501_3120 & ~v3_1517448501_3124;
   assign v3_1517448501_3127 = ~v3_1517448501_3128;
   assign v3_1517448501_3128 = ~v3_1517448501_1241 & ~v3_1517448501_3122;
   assign v3_1517448501_3129 = v3_1517448501_1251 & v3_1517448501_3127;
   assign v3_1517448501_3130 = ~v3_1517448501_3131;
   assign v3_1517448501_3131 = ~v3_1517448501_3125 & ~v3_1517448501_3129;
   assign v3_1517448501_3132 = ~v3_1517448501_3133;
   assign v3_1517448501_3133 = ~v3_1517448501_1251 & ~v3_1517448501_3127;
   assign v3_1517448501_3134 = v3_1517448501_1258 & v3_1517448501_3132;
   assign v3_1517448501_3135 = ~v3_1517448501_3136;
   assign v3_1517448501_3136 = ~v3_1517448501_3130 & ~v3_1517448501_3134;
   assign v3_1517448501_3137 = ~v3_1517448501_3138;
   assign v3_1517448501_3138 = ~v3_1517448501_1258 & ~v3_1517448501_3132;
   assign v3_1517448501_3139 = v3_1517448501_1263 & v3_1517448501_3137;
   assign v3_1517448501_3140 = ~v3_1517448501_3141;
   assign v3_1517448501_3141 = ~v3_1517448501_3135 & ~v3_1517448501_3139;
   assign v3_1517448501_3142 = v3_1517448501_3110 & ~v3_1517448501_3140;
   assign v3_1517448501_3143 = ~v3_1517448501_3144;
   assign v3_1517448501_3144 = ~v3_1517448501_1263 & ~v3_1517448501_3137;
   assign v3_1517448501_3145 = v3_1517448501_3142 & v3_1517448501_3143;
   assign v3_1517448501_3146 = v3_1517448501_2946 & v3_1517448501_3145;
   assign v3_1517448501_3147 = v3_1517448501_3146 & ~dve_invalid;
   assign v3_1517448501_3148 = 1'b0; 

   // Output Net Assignments
   assign id78 = v3_1517448501_80;

   // Property
   wire prop = !id78;
   wire prop_neg = !prop;
   assert property ( prop );

   // Non-blocking Assignments
   always @ (posedge v3_clock) begin
      v_m_initiator_0 <= v3_1517448501_139;
      v_party_nonce_initiator_0 <= v3_1517448501_170;
      v_m_initiator_1 <= v3_1517448501_183;
      v_party_nonce_initiator_1 <= v3_1517448501_213;
      v_m_initiator_2 <= v3_1517448501_226;
      v_party_nonce_initiator_2 <= v3_1517448501_256;
      v_m_responder_0 <= v3_1517448501_361;
      v_party_responder_0 <= v3_1517448501_391;
      v_party_nonce_responder_0 <= v3_1517448501_404;
      v_m_responder_1 <= v3_1517448501_461;
      v_party_responder_1 <= v3_1517448501_491;
      v_party_nonce_responder_1 <= v3_1517448501_504;
      v_m_responder_2 <= v3_1517448501_561;
      v_party_responder_2 <= v3_1517448501_591;
      v_party_nonce_responder_2 <= v3_1517448501_604;
      v_kNa <= v3_1517448501_610;
      v_kNb <= v3_1517448501_615;
      v_k_Na_Nb__A <= v3_1517448501_618;
      v_k_Na_A__B <= v3_1517448501_621;
      v_k_Nb__B <= v3_1517448501_626;
      v_m_intruder <= v3_1517448501_645;
      a_start_initiator_0 <= ~v3_1517448501_650;
      a_wait_resp_initiator_0 <= v3_1517448501_665;
      a_got_resp_initiator_0 <= v3_1517448501_680;
      a_commited_initiator_0 <= v3_1517448501_688;
      a_finished_initiator_0 <= v3_1517448501_696;
      a_corrupted_initiator_0 <= v3_1517448501_699;
      a_start_initiator_1 <= ~v3_1517448501_705;
      a_wait_resp_initiator_1 <= v3_1517448501_720;
      a_got_resp_initiator_1 <= v3_1517448501_735;
      a_commited_initiator_1 <= v3_1517448501_743;
      a_finished_initiator_1 <= v3_1517448501_751;
      a_corrupted_initiator_1 <= v3_1517448501_754;
      a_start_initiator_2 <= ~v3_1517448501_760;
      a_wait_resp_initiator_2 <= v3_1517448501_775;
      a_got_resp_initiator_2 <= v3_1517448501_790;
      a_commited_initiator_2 <= v3_1517448501_798;
      a_finished_initiator_2 <= v3_1517448501_806;
      a_corrupted_initiator_2 <= v3_1517448501_809;
      a_start_responder_0 <= ~v3_1517448501_835;
      a_got_msg_responder_0 <= v3_1517448501_886;
      a_send_reply_responder_0 <= v3_1517448501_894;
      a_wait_resp_responder_0 <= v3_1517448501_907;
      a_got_resp_responder_0 <= v3_1517448501_919;
      a_finished_responder_0 <= v3_1517448501_922;
      a_corrupted_responder_0 <= v3_1517448501_927;
      a_start_responder_1 <= ~v3_1517448501_953;
      a_got_msg_responder_1 <= v3_1517448501_1004;
      a_send_reply_responder_1 <= v3_1517448501_1012;
      a_wait_resp_responder_1 <= v3_1517448501_1025;
      a_got_resp_responder_1 <= v3_1517448501_1037;
      a_finished_responder_1 <= v3_1517448501_1040;
      a_corrupted_responder_1 <= v3_1517448501_1045;
      a_start_responder_2 <= ~v3_1517448501_1071;
      a_got_msg_responder_2 <= v3_1517448501_1122;
      a_send_reply_responder_2 <= v3_1517448501_1130;
      a_wait_resp_responder_2 <= v3_1517448501_1143;
      a_got_resp_responder_2 <= v3_1517448501_1155;
      a_finished_responder_2 <= v3_1517448501_1158;
      a_corrupted_responder_2 <= v3_1517448501_1163;
      a_q <= ~v3_1517448501_1201;
      a_got3 <= v3_1517448501_1218;
      a_c1 <= v3_1517448501_1226;
      a_c2 <= v3_1517448501_1235;
      a_d1 <= v3_1517448501_1241;
      a_got2 <= v3_1517448501_1251;
      a_e1 <= v3_1517448501_1258;
      a_f1 <= v3_1517448501_1263;
      dve_invalid <= ~v3_1517448501_3147;
   end
endmodule
