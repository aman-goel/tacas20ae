// RTL (Verilog) generated @ Wed Jan 31 20:28:21 2018 by V3 
//               compiled @ Jan 31 2018 12:00:50
// Internal nets are renamed with prefix "v3_1517448501_".

// Module needham
module needham
(
   v3_clock,
   f88,
   f86,
   f84,
   f81,
   f78,
   f00,
   f89,
   f87,
   f85,
   f82,
   f79,
   f02,
   f96,
   f93,
   f90,
   f76,
   f74,
   f72,
   f70,
   f68,
   f66,
   f64,
   f62,
   f60,
   f58,
   f56,
   f54,
   f52,
   f50,
   f48,
   f46,
   f44,
   f42,
   f40,
   f38,
   f36,
   f33,
   f30,
   f04,
   f97,
   f94,
   f91,
   f77,
   f75,
   f73,
   f71,
   f69,
   f67,
   f65,
   f63,
   f61,
   f59,
   f57,
   f55,
   f53,
   f51,
   f49,
   f47,
   f45,
   f43,
   f41,
   f39,
   f37,
   f34,
   f31,
   f08,
   f25,
   f15,
   f26,
   f16,
   f21,
   f20,
   f28,
   f18,
   f95,
   f92,
   f83,
   f80,
   f35,
   f32,
   f01,
   f03,
   f05,
   f06,
   f07,
   f09,
   f10,
   f11,
   f12,
   f19,
   f22,
   f27,
   f29,
   f13,
   f14,
   f17,
   f23,
   f24,
   id60
);

   // Clock Signal for Synchronous DFF
   input v3_clock;

   // I/O Declarations
   input f88;
   input f86;
   input f84;
   input f81;
   input f78;
   input f00;
   input f89;
   input f87;
   input f85;
   input f82;
   input f79;
   input f02;
   input f96;
   input f93;
   input f90;
   input f76;
   input f74;
   input f72;
   input f70;
   input f68;
   input f66;
   input f64;
   input f62;
   input f60;
   input f58;
   input f56;
   input f54;
   input f52;
   input f50;
   input f48;
   input f46;
   input f44;
   input f42;
   input f40;
   input f38;
   input f36;
   input f33;
   input f30;
   input f04;
   input f97;
   input f94;
   input f91;
   input f77;
   input f75;
   input f73;
   input f71;
   input f69;
   input f67;
   input f65;
   input f63;
   input f61;
   input f59;
   input f57;
   input f55;
   input f53;
   input f51;
   input f49;
   input f47;
   input f45;
   input f43;
   input f41;
   input f39;
   input f37;
   input f34;
   input f31;
   input f08;
   input f25;
   input f15;
   input f26;
   input f16;
   input f21;
   input f20;
   input f28;
   input f18;
   input f95;
   input f92;
   input f83;
   input f80;
   input f35;
   input f32;
   input f01;
   input f03;
   input f05;
   input f06;
   input f07;
   input f09;
   input f10;
   input f11;
   input f12;
   input f19;
   input f22;
   input f27;
   input f29;
   input f13;
   input f14;
   input f17;
   input f23;
   input f24;
   output id60;

   // Wire and Reg Declarations
   wire id0;
   reg [15:0] v_m_initiator_0 = 0;
   reg [15:0] v_party_nonce_initiator_0 = 0;
   reg [15:0] v_m_initiator_1 = 0;
   reg [15:0] v_party_nonce_initiator_1 = 0;
   reg [15:0] v_m_responder_0 = 0;
   reg [15:0] v_party_responder_0 = 0;
   reg [15:0] v_party_nonce_responder_0 = 0;
   reg [15:0] v_m_responder_1 = 0;
   reg [15:0] v_party_responder_1 = 0;
   reg [15:0] v_party_nonce_responder_1 = 0;
   reg [7:0] v_kNa = 0;
   reg [7:0] v_kNb = 0;
   reg [7:0] v_k_Na_Nb__A = 0;
   reg [7:0] v_k_Na_A__B = 0;
   reg [7:0] v_k_Nb__B = 0;
   reg [15:0] v_m_intruder = 0;
   reg a_start_initiator_0 = 0;
   reg a_wait_resp_initiator_0 = 0;
   reg a_got_resp_initiator_0 = 0;
   reg a_commited_initiator_0 = 0;
   reg a_finished_initiator_0 = 0;
   reg a_corrupted_initiator_0 = 0;
   reg a_start_initiator_1 = 0;
   reg a_wait_resp_initiator_1 = 0;
   reg a_got_resp_initiator_1 = 0;
   reg a_commited_initiator_1 = 0;
   reg a_finished_initiator_1 = 0;
   reg a_corrupted_initiator_1 = 0;
   reg a_start_responder_0 = 0;
   reg a_got_msg_responder_0 = 0;
   reg a_send_reply_responder_0 = 0;
   reg a_wait_resp_responder_0 = 0;
   reg a_got_resp_responder_0 = 0;
   reg a_finished_responder_0 = 0;
   reg a_corrupted_responder_0 = 0;
   reg a_start_responder_1 = 0;
   reg a_got_msg_responder_1 = 0;
   reg a_send_reply_responder_1 = 0;
   reg a_wait_resp_responder_1 = 0;
   reg a_got_resp_responder_1 = 0;
   reg a_finished_responder_1 = 0;
   reg a_corrupted_responder_1 = 0;
   reg a_q = 0;
   reg a_got3 = 0;
   reg a_c1 = 0;
   reg a_c2 = 0;
   reg a_d1 = 0;
   reg a_got2 = 0;
   reg a_e1 = 0;
   reg a_f1 = 0;
   reg dve_invalid = 0;
   wire [31:0] v3_1517448501_52;
   wire [15:0] v3_1517448501_53;
   wire [31:0] v3_1517448501_54;
   wire [4:0] v3_1517448501_55;
   wire [31:0] v3_1517448501_56;
   wire [31:0] v3_1517448501_57;
   wire [31:0] v3_1517448501_58;
   wire v3_1517448501_59;
   wire v3_1517448501_60;
   wire v3_1517448501_61;
   wire v3_1517448501_62;
   wire f88;
   wire [15:0] v3_1517448501_64;
   wire f86;
   wire [15:0] v3_1517448501_66;
   wire f84;
   wire [15:0] v3_1517448501_68;
   wire f81;
   wire [31:0] v3_1517448501_70;
   wire [31:0] v3_1517448501_71;
   wire [31:0] v3_1517448501_72;
   wire [31:0] v3_1517448501_73;
   wire [31:0] v3_1517448501_74;
   wire v3_1517448501_75;
   wire [31:0] v3_1517448501_76;
   wire [31:0] v3_1517448501_77;
   wire [31:0] v3_1517448501_78;
   wire [31:0] v3_1517448501_79;
   wire [31:0] v3_1517448501_80;
   wire [31:0] v3_1517448501_81;
   wire v3_1517448501_82;
   wire [31:0] v3_1517448501_83;
   wire [31:0] v3_1517448501_84;
   wire [31:0] v3_1517448501_85;
   wire [15:0] v3_1517448501_86;
   wire f78;
   wire [31:0] v3_1517448501_88;
   wire [31:0] v3_1517448501_89;
   wire [31:0] v3_1517448501_90;
   wire [31:0] v3_1517448501_91;
   wire [31:0] v3_1517448501_92;
   wire v3_1517448501_93;
   wire [31:0] v3_1517448501_94;
   wire [31:0] v3_1517448501_95;
   wire [31:0] v3_1517448501_96;
   wire [31:0] v3_1517448501_97;
   wire [15:0] v3_1517448501_98;
   wire [15:0] v3_1517448501_99;
   wire [15:0] v3_1517448501_100;
   wire [15:0] v3_1517448501_101;
   wire [15:0] v3_1517448501_102;
   wire [15:0] v3_1517448501_103;
   wire [15:0] v3_1517448501_104;
   wire f00;
   wire [31:0] v3_1517448501_106;
   wire [31:0] v3_1517448501_107;
   wire [31:0] v3_1517448501_108;
   wire [31:0] v3_1517448501_109;
   wire v3_1517448501_110;
   wire [31:0] v3_1517448501_111;
   wire [31:0] v3_1517448501_112;
   wire v3_1517448501_113;
   wire v3_1517448501_114;
   wire [31:0] v3_1517448501_115;
   wire [31:0] v3_1517448501_116;
   wire [31:0] v3_1517448501_117;
   wire [31:0] v3_1517448501_118;
   wire [31:0] v3_1517448501_119;
   wire [31:0] v3_1517448501_120;
   wire [31:0] v3_1517448501_121;
   wire [31:0] v3_1517448501_122;
   wire v3_1517448501_123;
   wire v3_1517448501_124;
   wire v3_1517448501_125;
   wire [31:0] v3_1517448501_126;
   wire [31:0] v3_1517448501_127;
   wire [31:0] v3_1517448501_128;
   wire [31:0] v3_1517448501_129;
   wire [31:0] v3_1517448501_130;
   wire [31:0] v3_1517448501_131;
   wire [31:0] v3_1517448501_132;
   wire [15:0] v3_1517448501_133;
   wire [15:0] v3_1517448501_134;
   wire [15:0] v3_1517448501_135;
   wire f89;
   wire f87;
   wire f85;
   wire f82;
   wire f79;
   wire [15:0] v3_1517448501_141;
   wire [15:0] v3_1517448501_142;
   wire [15:0] v3_1517448501_143;
   wire [15:0] v3_1517448501_144;
   wire [15:0] v3_1517448501_145;
   wire [15:0] v3_1517448501_146;
   wire f02;
   wire [31:0] v3_1517448501_148;
   wire [31:0] v3_1517448501_149;
   wire [31:0] v3_1517448501_150;
   wire [31:0] v3_1517448501_151;
   wire v3_1517448501_152;
   wire [31:0] v3_1517448501_153;
   wire v3_1517448501_154;
   wire v3_1517448501_155;
   wire [31:0] v3_1517448501_156;
   wire [31:0] v3_1517448501_157;
   wire [31:0] v3_1517448501_158;
   wire [31:0] v3_1517448501_159;
   wire [31:0] v3_1517448501_160;
   wire [31:0] v3_1517448501_161;
   wire [31:0] v3_1517448501_162;
   wire [31:0] v3_1517448501_163;
   wire v3_1517448501_164;
   wire v3_1517448501_165;
   wire v3_1517448501_166;
   wire [31:0] v3_1517448501_167;
   wire [31:0] v3_1517448501_168;
   wire [31:0] v3_1517448501_169;
   wire [31:0] v3_1517448501_170;
   wire [31:0] v3_1517448501_171;
   wire [31:0] v3_1517448501_172;
   wire [31:0] v3_1517448501_173;
   wire [15:0] v3_1517448501_174;
   wire [15:0] v3_1517448501_175;
   wire [15:0] v3_1517448501_176;
   wire f96;
   wire [15:0] v3_1517448501_178;
   wire f93;
   wire [31:0] v3_1517448501_180;
   wire [31:0] v3_1517448501_181;
   wire [31:0] v3_1517448501_182;
   wire [31:0] v3_1517448501_183;
   wire [31:0] v3_1517448501_184;
   wire v3_1517448501_185;
   wire [31:0] v3_1517448501_186;
   wire [15:0] v3_1517448501_187;
   wire f90;
   wire [31:0] v3_1517448501_189;
   wire [31:0] v3_1517448501_190;
   wire [31:0] v3_1517448501_191;
   wire [31:0] v3_1517448501_192;
   wire [31:0] v3_1517448501_193;
   wire v3_1517448501_194;
   wire [31:0] v3_1517448501_195;
   wire [15:0] v3_1517448501_196;
   wire f76;
   wire [15:0] v3_1517448501_198;
   wire f74;
   wire [15:0] v3_1517448501_200;
   wire f72;
   wire [15:0] v3_1517448501_202;
   wire f70;
   wire [15:0] v3_1517448501_204;
   wire f68;
   wire [15:0] v3_1517448501_206;
   wire f66;
   wire [15:0] v3_1517448501_208;
   wire f64;
   wire [15:0] v3_1517448501_210;
   wire f62;
   wire [15:0] v3_1517448501_212;
   wire f60;
   wire [15:0] v3_1517448501_214;
   wire f58;
   wire [15:0] v3_1517448501_216;
   wire f56;
   wire [15:0] v3_1517448501_218;
   wire f54;
   wire [15:0] v3_1517448501_220;
   wire f52;
   wire [15:0] v3_1517448501_222;
   wire f50;
   wire [15:0] v3_1517448501_224;
   wire f48;
   wire [15:0] v3_1517448501_226;
   wire f46;
   wire [15:0] v3_1517448501_228;
   wire f44;
   wire [15:0] v3_1517448501_230;
   wire f42;
   wire [15:0] v3_1517448501_232;
   wire f40;
   wire [15:0] v3_1517448501_234;
   wire f38;
   wire [15:0] v3_1517448501_236;
   wire f36;
   wire [15:0] v3_1517448501_238;
   wire f33;
   wire [15:0] v3_1517448501_240;
   wire f30;
   wire [15:0] v3_1517448501_242;
   wire [15:0] v3_1517448501_243;
   wire [15:0] v3_1517448501_244;
   wire [15:0] v3_1517448501_245;
   wire [15:0] v3_1517448501_246;
   wire [15:0] v3_1517448501_247;
   wire [15:0] v3_1517448501_248;
   wire [15:0] v3_1517448501_249;
   wire [15:0] v3_1517448501_250;
   wire [15:0] v3_1517448501_251;
   wire [15:0] v3_1517448501_252;
   wire [15:0] v3_1517448501_253;
   wire [15:0] v3_1517448501_254;
   wire [15:0] v3_1517448501_255;
   wire [15:0] v3_1517448501_256;
   wire [15:0] v3_1517448501_257;
   wire [15:0] v3_1517448501_258;
   wire [15:0] v3_1517448501_259;
   wire [15:0] v3_1517448501_260;
   wire [15:0] v3_1517448501_261;
   wire [15:0] v3_1517448501_262;
   wire [15:0] v3_1517448501_263;
   wire [15:0] v3_1517448501_264;
   wire [15:0] v3_1517448501_265;
   wire [15:0] v3_1517448501_266;
   wire [15:0] v3_1517448501_267;
   wire [15:0] v3_1517448501_268;
   wire f04;
   wire [31:0] v3_1517448501_270;
   wire [31:0] v3_1517448501_271;
   wire [31:0] v3_1517448501_272;
   wire [31:0] v3_1517448501_273;
   wire v3_1517448501_274;
   wire [31:0] v3_1517448501_275;
   wire v3_1517448501_276;
   wire v3_1517448501_277;
   wire [31:0] v3_1517448501_278;
   wire [31:0] v3_1517448501_279;
   wire [31:0] v3_1517448501_280;
   wire [31:0] v3_1517448501_281;
   wire [31:0] v3_1517448501_282;
   wire [31:0] v3_1517448501_283;
   wire [31:0] v3_1517448501_284;
   wire [31:0] v3_1517448501_285;
   wire v3_1517448501_286;
   wire v3_1517448501_287;
   wire v3_1517448501_288;
   wire [31:0] v3_1517448501_289;
   wire [31:0] v3_1517448501_290;
   wire [31:0] v3_1517448501_291;
   wire [31:0] v3_1517448501_292;
   wire [31:0] v3_1517448501_293;
   wire [31:0] v3_1517448501_294;
   wire [31:0] v3_1517448501_295;
   wire [15:0] v3_1517448501_296;
   wire [15:0] v3_1517448501_297;
   wire [15:0] v3_1517448501_298;
   wire [31:0] v3_1517448501_299;
   wire v3_1517448501_300;
   wire v3_1517448501_301;
   wire [31:0] v3_1517448501_302;
   wire [31:0] v3_1517448501_303;
   wire [31:0] v3_1517448501_304;
   wire [31:0] v3_1517448501_305;
   wire [31:0] v3_1517448501_306;
   wire [31:0] v3_1517448501_307;
   wire [31:0] v3_1517448501_308;
   wire [15:0] v3_1517448501_309;
   wire [15:0] v3_1517448501_310;
   wire [15:0] v3_1517448501_311;
   wire f97;
   wire f94;
   wire f91;
   wire f77;
   wire f75;
   wire f73;
   wire f71;
   wire f69;
   wire f67;
   wire f65;
   wire f63;
   wire f61;
   wire f59;
   wire f57;
   wire f55;
   wire f53;
   wire f51;
   wire f49;
   wire f47;
   wire f45;
   wire f43;
   wire f41;
   wire f39;
   wire f37;
   wire f34;
   wire f31;
   wire [15:0] v3_1517448501_338;
   wire [15:0] v3_1517448501_339;
   wire [15:0] v3_1517448501_340;
   wire [15:0] v3_1517448501_341;
   wire [15:0] v3_1517448501_342;
   wire [15:0] v3_1517448501_343;
   wire [15:0] v3_1517448501_344;
   wire [15:0] v3_1517448501_345;
   wire [15:0] v3_1517448501_346;
   wire [15:0] v3_1517448501_347;
   wire [15:0] v3_1517448501_348;
   wire [15:0] v3_1517448501_349;
   wire [15:0] v3_1517448501_350;
   wire [15:0] v3_1517448501_351;
   wire [15:0] v3_1517448501_352;
   wire [15:0] v3_1517448501_353;
   wire [15:0] v3_1517448501_354;
   wire [15:0] v3_1517448501_355;
   wire [15:0] v3_1517448501_356;
   wire [15:0] v3_1517448501_357;
   wire [15:0] v3_1517448501_358;
   wire [15:0] v3_1517448501_359;
   wire [15:0] v3_1517448501_360;
   wire [15:0] v3_1517448501_361;
   wire [15:0] v3_1517448501_362;
   wire [15:0] v3_1517448501_363;
   wire [15:0] v3_1517448501_364;
   wire f08;
   wire [31:0] v3_1517448501_366;
   wire [31:0] v3_1517448501_367;
   wire [31:0] v3_1517448501_368;
   wire [31:0] v3_1517448501_369;
   wire v3_1517448501_370;
   wire [31:0] v3_1517448501_371;
   wire v3_1517448501_372;
   wire v3_1517448501_373;
   wire [31:0] v3_1517448501_374;
   wire [31:0] v3_1517448501_375;
   wire [31:0] v3_1517448501_376;
   wire [31:0] v3_1517448501_377;
   wire [31:0] v3_1517448501_378;
   wire [31:0] v3_1517448501_379;
   wire [31:0] v3_1517448501_380;
   wire [31:0] v3_1517448501_381;
   wire v3_1517448501_382;
   wire v3_1517448501_383;
   wire v3_1517448501_384;
   wire [31:0] v3_1517448501_385;
   wire [31:0] v3_1517448501_386;
   wire [31:0] v3_1517448501_387;
   wire [31:0] v3_1517448501_388;
   wire [31:0] v3_1517448501_389;
   wire [31:0] v3_1517448501_390;
   wire [31:0] v3_1517448501_391;
   wire [15:0] v3_1517448501_392;
   wire [15:0] v3_1517448501_393;
   wire [15:0] v3_1517448501_394;
   wire [31:0] v3_1517448501_395;
   wire v3_1517448501_396;
   wire v3_1517448501_397;
   wire [31:0] v3_1517448501_398;
   wire [31:0] v3_1517448501_399;
   wire [31:0] v3_1517448501_400;
   wire [31:0] v3_1517448501_401;
   wire [31:0] v3_1517448501_402;
   wire [31:0] v3_1517448501_403;
   wire [31:0] v3_1517448501_404;
   wire [15:0] v3_1517448501_405;
   wire [15:0] v3_1517448501_406;
   wire [15:0] v3_1517448501_407;
   wire f25;
   wire [7:0] v3_1517448501_409;
   wire f15;
   wire [7:0] v3_1517448501_411;
   wire [7:0] v3_1517448501_412;
   wire [7:0] v3_1517448501_413;
   wire f26;
   wire f16;
   wire [7:0] v3_1517448501_416;
   wire [7:0] v3_1517448501_417;
   wire [7:0] v3_1517448501_418;
   wire f21;
   wire [7:0] v3_1517448501_420;
   wire [7:0] v3_1517448501_421;
   wire f20;
   wire [7:0] v3_1517448501_423;
   wire [7:0] v3_1517448501_424;
   wire f28;
   wire f18;
   wire [7:0] v3_1517448501_427;
   wire [7:0] v3_1517448501_428;
   wire [7:0] v3_1517448501_429;
   wire f95;
   wire f92;
   wire f83;
   wire f80;
   wire f35;
   wire f32;
   wire [15:0] v3_1517448501_436;
   wire [15:0] v3_1517448501_437;
   wire [15:0] v3_1517448501_438;
   wire [15:0] v3_1517448501_439;
   wire [15:0] v3_1517448501_440;
   wire [15:0] v3_1517448501_441;
   wire [15:0] v3_1517448501_442;
   wire v3_1517448501_443;
   wire v3_1517448501_444;
   wire v3_1517448501_445;
   wire v3_1517448501_446;
   wire v3_1517448501_447;
   wire v3_1517448501_448;
   wire v3_1517448501_449;
   wire v3_1517448501_450;
   wire v3_1517448501_451;
   wire v3_1517448501_452;
   wire v3_1517448501_453;
   wire v3_1517448501_454;
   wire v3_1517448501_455;
   wire v3_1517448501_456;
   wire v3_1517448501_457;
   wire v3_1517448501_458;
   wire v3_1517448501_459;
   wire f01;
   wire v3_1517448501_461;
   wire v3_1517448501_462;
   wire v3_1517448501_463;
   wire v3_1517448501_464;
   wire v3_1517448501_465;
   wire v3_1517448501_466;
   wire v3_1517448501_467;
   wire v3_1517448501_468;
   wire v3_1517448501_469;
   wire v3_1517448501_470;
   wire v3_1517448501_471;
   wire v3_1517448501_472;
   wire v3_1517448501_473;
   wire v3_1517448501_474;
   wire v3_1517448501_475;
   wire v3_1517448501_476;
   wire v3_1517448501_477;
   wire v3_1517448501_478;
   wire v3_1517448501_479;
   wire v3_1517448501_480;
   wire v3_1517448501_481;
   wire v3_1517448501_482;
   wire v3_1517448501_483;
   wire v3_1517448501_484;
   wire v3_1517448501_485;
   wire v3_1517448501_486;
   wire v3_1517448501_487;
   wire v3_1517448501_488;
   wire v3_1517448501_489;
   wire v3_1517448501_490;
   wire v3_1517448501_491;
   wire v3_1517448501_492;
   wire v3_1517448501_493;
   wire v3_1517448501_494;
   wire v3_1517448501_495;
   wire v3_1517448501_496;
   wire v3_1517448501_497;
   wire v3_1517448501_498;
   wire v3_1517448501_499;
   wire v3_1517448501_500;
   wire v3_1517448501_501;
   wire v3_1517448501_502;
   wire v3_1517448501_503;
   wire v3_1517448501_504;
   wire v3_1517448501_505;
   wire f03;
   wire v3_1517448501_507;
   wire v3_1517448501_508;
   wire v3_1517448501_509;
   wire v3_1517448501_510;
   wire v3_1517448501_511;
   wire v3_1517448501_512;
   wire v3_1517448501_513;
   wire v3_1517448501_514;
   wire v3_1517448501_515;
   wire v3_1517448501_516;
   wire v3_1517448501_517;
   wire v3_1517448501_518;
   wire v3_1517448501_519;
   wire v3_1517448501_520;
   wire v3_1517448501_521;
   wire v3_1517448501_522;
   wire v3_1517448501_523;
   wire v3_1517448501_524;
   wire v3_1517448501_525;
   wire v3_1517448501_526;
   wire v3_1517448501_527;
   wire v3_1517448501_528;
   wire v3_1517448501_529;
   wire v3_1517448501_530;
   wire v3_1517448501_531;
   wire v3_1517448501_532;
   wire v3_1517448501_533;
   wire v3_1517448501_534;
   wire v3_1517448501_535;
   wire v3_1517448501_536;
   wire v3_1517448501_537;
   wire v3_1517448501_538;
   wire v3_1517448501_539;
   wire v3_1517448501_540;
   wire v3_1517448501_541;
   wire v3_1517448501_542;
   wire v3_1517448501_543;
   wire v3_1517448501_544;
   wire v3_1517448501_545;
   wire v3_1517448501_546;
   wire v3_1517448501_547;
   wire v3_1517448501_548;
   wire v3_1517448501_549;
   wire v3_1517448501_550;
   wire v3_1517448501_551;
   wire v3_1517448501_552;
   wire v3_1517448501_553;
   wire v3_1517448501_554;
   wire v3_1517448501_555;
   wire v3_1517448501_556;
   wire v3_1517448501_557;
   wire v3_1517448501_558;
   wire v3_1517448501_559;
   wire f05;
   wire v3_1517448501_561;
   wire v3_1517448501_562;
   wire v3_1517448501_563;
   wire v3_1517448501_564;
   wire v3_1517448501_565;
   wire v3_1517448501_566;
   wire v3_1517448501_567;
   wire v3_1517448501_568;
   wire v3_1517448501_569;
   wire v3_1517448501_570;
   wire v3_1517448501_571;
   wire v3_1517448501_572;
   wire v3_1517448501_573;
   wire v3_1517448501_574;
   wire v3_1517448501_575;
   wire v3_1517448501_576;
   wire v3_1517448501_577;
   wire v3_1517448501_578;
   wire v3_1517448501_579;
   wire v3_1517448501_580;
   wire v3_1517448501_581;
   wire v3_1517448501_582;
   wire v3_1517448501_583;
   wire v3_1517448501_584;
   wire v3_1517448501_585;
   wire v3_1517448501_586;
   wire v3_1517448501_587;
   wire v3_1517448501_588;
   wire v3_1517448501_589;
   wire v3_1517448501_590;
   wire v3_1517448501_591;
   wire v3_1517448501_592;
   wire v3_1517448501_593;
   wire v3_1517448501_594;
   wire v3_1517448501_595;
   wire v3_1517448501_596;
   wire v3_1517448501_597;
   wire v3_1517448501_598;
   wire v3_1517448501_599;
   wire v3_1517448501_600;
   wire v3_1517448501_601;
   wire v3_1517448501_602;
   wire v3_1517448501_603;
   wire v3_1517448501_604;
   wire v3_1517448501_605;
   wire v3_1517448501_606;
   wire v3_1517448501_607;
   wire v3_1517448501_608;
   wire v3_1517448501_609;
   wire v3_1517448501_610;
   wire v3_1517448501_611;
   wire v3_1517448501_612;
   wire v3_1517448501_613;
   wire v3_1517448501_614;
   wire v3_1517448501_615;
   wire v3_1517448501_616;
   wire v3_1517448501_617;
   wire v3_1517448501_618;
   wire v3_1517448501_619;
   wire v3_1517448501_620;
   wire v3_1517448501_621;
   wire v3_1517448501_622;
   wire v3_1517448501_623;
   wire v3_1517448501_624;
   wire f06;
   wire v3_1517448501_626;
   wire f07;
   wire v3_1517448501_628;
   wire v3_1517448501_629;
   wire v3_1517448501_630;
   wire v3_1517448501_631;
   wire v3_1517448501_632;
   wire v3_1517448501_633;
   wire v3_1517448501_634;
   wire v3_1517448501_635;
   wire v3_1517448501_636;
   wire v3_1517448501_637;
   wire v3_1517448501_638;
   wire v3_1517448501_639;
   wire v3_1517448501_640;
   wire v3_1517448501_641;
   wire v3_1517448501_642;
   wire v3_1517448501_643;
   wire v3_1517448501_644;
   wire v3_1517448501_645;
   wire v3_1517448501_646;
   wire v3_1517448501_647;
   wire v3_1517448501_648;
   wire v3_1517448501_649;
   wire v3_1517448501_650;
   wire v3_1517448501_651;
   wire v3_1517448501_652;
   wire v3_1517448501_653;
   wire v3_1517448501_654;
   wire v3_1517448501_655;
   wire v3_1517448501_656;
   wire v3_1517448501_657;
   wire v3_1517448501_658;
   wire v3_1517448501_659;
   wire v3_1517448501_660;
   wire v3_1517448501_661;
   wire v3_1517448501_662;
   wire v3_1517448501_663;
   wire v3_1517448501_664;
   wire v3_1517448501_665;
   wire v3_1517448501_666;
   wire v3_1517448501_667;
   wire v3_1517448501_668;
   wire f09;
   wire v3_1517448501_670;
   wire v3_1517448501_671;
   wire v3_1517448501_672;
   wire v3_1517448501_673;
   wire v3_1517448501_674;
   wire v3_1517448501_675;
   wire v3_1517448501_676;
   wire v3_1517448501_677;
   wire v3_1517448501_678;
   wire v3_1517448501_679;
   wire v3_1517448501_680;
   wire v3_1517448501_681;
   wire v3_1517448501_682;
   wire v3_1517448501_683;
   wire v3_1517448501_684;
   wire v3_1517448501_685;
   wire v3_1517448501_686;
   wire v3_1517448501_687;
   wire v3_1517448501_688;
   wire v3_1517448501_689;
   wire v3_1517448501_690;
   wire v3_1517448501_691;
   wire v3_1517448501_692;
   wire v3_1517448501_693;
   wire v3_1517448501_694;
   wire v3_1517448501_695;
   wire v3_1517448501_696;
   wire v3_1517448501_697;
   wire v3_1517448501_698;
   wire v3_1517448501_699;
   wire v3_1517448501_700;
   wire v3_1517448501_701;
   wire v3_1517448501_702;
   wire v3_1517448501_703;
   wire v3_1517448501_704;
   wire v3_1517448501_705;
   wire v3_1517448501_706;
   wire v3_1517448501_707;
   wire v3_1517448501_708;
   wire v3_1517448501_709;
   wire v3_1517448501_710;
   wire v3_1517448501_711;
   wire v3_1517448501_712;
   wire v3_1517448501_713;
   wire v3_1517448501_714;
   wire v3_1517448501_715;
   wire v3_1517448501_716;
   wire v3_1517448501_717;
   wire v3_1517448501_718;
   wire v3_1517448501_719;
   wire v3_1517448501_720;
   wire v3_1517448501_721;
   wire v3_1517448501_722;
   wire v3_1517448501_723;
   wire v3_1517448501_724;
   wire v3_1517448501_725;
   wire v3_1517448501_726;
   wire v3_1517448501_727;
   wire v3_1517448501_728;
   wire v3_1517448501_729;
   wire v3_1517448501_730;
   wire v3_1517448501_731;
   wire v3_1517448501_732;
   wire v3_1517448501_733;
   wire f10;
   wire v3_1517448501_735;
   wire f11;
   wire v3_1517448501_737;
   wire v3_1517448501_738;
   wire v3_1517448501_739;
   wire v3_1517448501_740;
   wire v3_1517448501_741;
   wire v3_1517448501_742;
   wire v3_1517448501_743;
   wire v3_1517448501_744;
   wire v3_1517448501_745;
   wire v3_1517448501_746;
   wire v3_1517448501_747;
   wire v3_1517448501_748;
   wire v3_1517448501_749;
   wire v3_1517448501_750;
   wire v3_1517448501_751;
   wire v3_1517448501_752;
   wire f12;
   wire v3_1517448501_754;
   wire v3_1517448501_755;
   wire v3_1517448501_756;
   wire v3_1517448501_757;
   wire f19;
   wire v3_1517448501_759;
   wire v3_1517448501_760;
   wire v3_1517448501_761;
   wire v3_1517448501_762;
   wire v3_1517448501_763;
   wire v3_1517448501_764;
   wire f22;
   wire v3_1517448501_766;
   wire v3_1517448501_767;
   wire v3_1517448501_768;
   wire v3_1517448501_769;
   wire v3_1517448501_770;
   wire v3_1517448501_771;
   wire f27;
   wire v3_1517448501_773;
   wire v3_1517448501_774;
   wire v3_1517448501_775;
   wire v3_1517448501_776;
   wire f29;
   wire v3_1517448501_778;
   wire v3_1517448501_779;
   wire v3_1517448501_780;
   wire v3_1517448501_781;
   wire v3_1517448501_782;
   wire v3_1517448501_783;
   wire v3_1517448501_784;
   wire v3_1517448501_785;
   wire v3_1517448501_786;
   wire v3_1517448501_787;
   wire f13;
   wire v3_1517448501_789;
   wire f14;
   wire v3_1517448501_791;
   wire v3_1517448501_792;
   wire v3_1517448501_793;
   wire v3_1517448501_794;
   wire v3_1517448501_795;
   wire v3_1517448501_796;
   wire v3_1517448501_797;
   wire v3_1517448501_798;
   wire v3_1517448501_799;
   wire v3_1517448501_800;
   wire v3_1517448501_801;
   wire v3_1517448501_802;
   wire v3_1517448501_803;
   wire v3_1517448501_804;
   wire f17;
   wire v3_1517448501_806;
   wire v3_1517448501_807;
   wire v3_1517448501_808;
   wire v3_1517448501_809;
   wire v3_1517448501_810;
   wire v3_1517448501_811;
   wire v3_1517448501_812;
   wire v3_1517448501_813;
   wire v3_1517448501_814;
   wire v3_1517448501_815;
   wire v3_1517448501_816;
   wire v3_1517448501_817;
   wire v3_1517448501_818;
   wire v3_1517448501_819;
   wire v3_1517448501_820;
   wire v3_1517448501_821;
   wire v3_1517448501_822;
   wire f23;
   wire v3_1517448501_824;
   wire f24;
   wire v3_1517448501_826;
   wire v3_1517448501_827;
   wire v3_1517448501_828;
   wire v3_1517448501_829;
   wire v3_1517448501_830;
   wire v3_1517448501_831;
   wire v3_1517448501_832;
   wire v3_1517448501_833;
   wire v3_1517448501_834;
   wire v3_1517448501_835;
   wire v3_1517448501_836;
   wire v3_1517448501_837;
   wire v3_1517448501_838;
   wire v3_1517448501_839;
   wire v3_1517448501_840;
   wire v3_1517448501_841;
   wire v3_1517448501_842;
   wire [31:0] v3_1517448501_843;
   wire [31:0] v3_1517448501_844;
   wire v3_1517448501_845;
   wire v3_1517448501_846;
   wire [31:0] v3_1517448501_847;
   wire [31:0] v3_1517448501_848;
   wire [31:0] v3_1517448501_849;
   wire [31:0] v3_1517448501_850;
   wire [31:0] v3_1517448501_851;
   wire [31:0] v3_1517448501_852;
   wire [31:0] v3_1517448501_853;
   wire v3_1517448501_854;
   wire [31:0] v3_1517448501_855;
   wire v3_1517448501_856;
   wire v3_1517448501_857;
   wire v3_1517448501_858;
   wire [31:0] v3_1517448501_859;
   wire [31:0] v3_1517448501_860;
   wire [31:0] v3_1517448501_861;
   wire [31:0] v3_1517448501_862;
   wire [31:0] v3_1517448501_863;
   wire [31:0] v3_1517448501_864;
   wire [31:0] v3_1517448501_865;
   wire v3_1517448501_866;
   wire v3_1517448501_867;
   wire v3_1517448501_868;
   wire v3_1517448501_869;
   wire v3_1517448501_870;
   wire v3_1517448501_871;
   wire v3_1517448501_872;
   wire v3_1517448501_873;
   wire v3_1517448501_874;
   wire [31:0] v3_1517448501_875;
   wire [31:0] v3_1517448501_876;
   wire v3_1517448501_877;
   wire v3_1517448501_878;
   wire [31:0] v3_1517448501_879;
   wire [31:0] v3_1517448501_880;
   wire [31:0] v3_1517448501_881;
   wire [31:0] v3_1517448501_882;
   wire [31:0] v3_1517448501_883;
   wire [31:0] v3_1517448501_884;
   wire [31:0] v3_1517448501_885;
   wire v3_1517448501_886;
   wire [31:0] v3_1517448501_887;
   wire [31:0] v3_1517448501_888;
   wire v3_1517448501_889;
   wire v3_1517448501_890;
   wire v3_1517448501_891;
   wire [31:0] v3_1517448501_892;
   wire [31:0] v3_1517448501_893;
   wire [31:0] v3_1517448501_894;
   wire [31:0] v3_1517448501_895;
   wire [31:0] v3_1517448501_896;
   wire [31:0] v3_1517448501_897;
   wire [31:0] v3_1517448501_898;
   wire v3_1517448501_899;
   wire v3_1517448501_900;
   wire v3_1517448501_901;
   wire v3_1517448501_902;
   wire v3_1517448501_903;
   wire v3_1517448501_904;
   wire v3_1517448501_905;
   wire v3_1517448501_906;
   wire v3_1517448501_907;
   wire v3_1517448501_908;
   wire [31:0] v3_1517448501_909;
   wire [31:0] v3_1517448501_910;
   wire v3_1517448501_911;
   wire v3_1517448501_912;
   wire v3_1517448501_913;
   wire [31:0] v3_1517448501_914;
   wire [31:0] v3_1517448501_915;
   wire [31:0] v3_1517448501_916;
   wire [31:0] v3_1517448501_917;
   wire [31:0] v3_1517448501_918;
   wire [31:0] v3_1517448501_919;
   wire [31:0] v3_1517448501_920;
   wire v3_1517448501_921;
   wire v3_1517448501_922;
   wire v3_1517448501_923;
   wire v3_1517448501_924;
   wire v3_1517448501_925;
   wire v3_1517448501_926;
   wire v3_1517448501_927;
   wire v3_1517448501_928;
   wire v3_1517448501_929;
   wire [31:0] v3_1517448501_930;
   wire v3_1517448501_931;
   wire v3_1517448501_932;
   wire v3_1517448501_933;
   wire v3_1517448501_934;
   wire v3_1517448501_935;
   wire v3_1517448501_936;
   wire v3_1517448501_937;
   wire v3_1517448501_938;
   wire v3_1517448501_939;
   wire v3_1517448501_940;
   wire v3_1517448501_941;
   wire [31:0] v3_1517448501_942;
   wire [31:0] v3_1517448501_943;
   wire v3_1517448501_944;
   wire v3_1517448501_945;
   wire v3_1517448501_946;
   wire [31:0] v3_1517448501_947;
   wire [31:0] v3_1517448501_948;
   wire [31:0] v3_1517448501_949;
   wire [31:0] v3_1517448501_950;
   wire [31:0] v3_1517448501_951;
   wire [31:0] v3_1517448501_952;
   wire [31:0] v3_1517448501_953;
   wire v3_1517448501_954;
   wire v3_1517448501_955;
   wire v3_1517448501_956;
   wire v3_1517448501_957;
   wire v3_1517448501_958;
   wire v3_1517448501_959;
   wire v3_1517448501_960;
   wire v3_1517448501_961;
   wire v3_1517448501_962;
   wire [31:0] v3_1517448501_963;
   wire v3_1517448501_964;
   wire v3_1517448501_965;
   wire v3_1517448501_966;
   wire v3_1517448501_967;
   wire v3_1517448501_968;
   wire v3_1517448501_969;
   wire v3_1517448501_970;
   wire v3_1517448501_971;
   wire v3_1517448501_972;
   wire v3_1517448501_973;
   wire v3_1517448501_974;
   wire v3_1517448501_975;
   wire v3_1517448501_976;
   wire v3_1517448501_977;
   wire [31:0] v3_1517448501_978;
   wire [31:0] v3_1517448501_979;
   wire [31:0] v3_1517448501_980;
   wire [31:0] v3_1517448501_981;
   wire v3_1517448501_982;
   wire [31:0] v3_1517448501_983;
   wire v3_1517448501_984;
   wire v3_1517448501_985;
   wire v3_1517448501_986;
   wire [31:0] v3_1517448501_987;
   wire [31:0] v3_1517448501_988;
   wire [31:0] v3_1517448501_989;
   wire [31:0] v3_1517448501_990;
   wire [31:0] v3_1517448501_991;
   wire [31:0] v3_1517448501_992;
   wire [31:0] v3_1517448501_993;
   wire v3_1517448501_994;
   wire v3_1517448501_995;
   wire v3_1517448501_996;
   wire v3_1517448501_997;
   wire v3_1517448501_998;
   wire v3_1517448501_999;
   wire v3_1517448501_1000;
   wire v3_1517448501_1001;
   wire v3_1517448501_1002;
   wire [31:0] v3_1517448501_1003;
   wire v3_1517448501_1004;
   wire v3_1517448501_1005;
   wire [31:0] v3_1517448501_1006;
   wire [31:0] v3_1517448501_1007;
   wire [31:0] v3_1517448501_1008;
   wire [31:0] v3_1517448501_1009;
   wire [31:0] v3_1517448501_1010;
   wire [31:0] v3_1517448501_1011;
   wire [31:0] v3_1517448501_1012;
   wire v3_1517448501_1013;
   wire v3_1517448501_1014;
   wire v3_1517448501_1015;
   wire v3_1517448501_1016;
   wire v3_1517448501_1017;
   wire v3_1517448501_1018;
   wire v3_1517448501_1019;
   wire v3_1517448501_1020;
   wire v3_1517448501_1021;
   wire v3_1517448501_1022;
   wire v3_1517448501_1023;
   wire v3_1517448501_1024;
   wire v3_1517448501_1025;
   wire v3_1517448501_1026;
   wire v3_1517448501_1027;
   wire [31:0] v3_1517448501_1028;
   wire v3_1517448501_1029;
   wire v3_1517448501_1030;
   wire [31:0] v3_1517448501_1031;
   wire [31:0] v3_1517448501_1032;
   wire [31:0] v3_1517448501_1033;
   wire [31:0] v3_1517448501_1034;
   wire [31:0] v3_1517448501_1035;
   wire [31:0] v3_1517448501_1036;
   wire [31:0] v3_1517448501_1037;
   wire [31:0] v3_1517448501_1038;
   wire v3_1517448501_1039;
   wire v3_1517448501_1040;
   wire v3_1517448501_1041;
   wire [31:0] v3_1517448501_1042;
   wire [31:0] v3_1517448501_1043;
   wire [31:0] v3_1517448501_1044;
   wire [31:0] v3_1517448501_1045;
   wire [31:0] v3_1517448501_1046;
   wire [31:0] v3_1517448501_1047;
   wire [31:0] v3_1517448501_1048;
   wire v3_1517448501_1049;
   wire v3_1517448501_1050;
   wire v3_1517448501_1051;
   wire v3_1517448501_1052;
   wire v3_1517448501_1053;
   wire v3_1517448501_1054;
   wire v3_1517448501_1055;
   wire v3_1517448501_1056;
   wire v3_1517448501_1057;
   wire v3_1517448501_1058;
   wire v3_1517448501_1059;
   wire v3_1517448501_1060;
   wire v3_1517448501_1061;
   wire v3_1517448501_1062;
   wire v3_1517448501_1063;
   wire v3_1517448501_1064;
   wire v3_1517448501_1065;
   wire v3_1517448501_1066;
   wire v3_1517448501_1067;
   wire v3_1517448501_1068;
   wire v3_1517448501_1069;
   wire v3_1517448501_1070;
   wire v3_1517448501_1071;
   wire v3_1517448501_1072;
   wire v3_1517448501_1073;
   wire v3_1517448501_1074;
   wire v3_1517448501_1075;
   wire v3_1517448501_1076;
   wire v3_1517448501_1077;
   wire v3_1517448501_1078;
   wire v3_1517448501_1079;
   wire v3_1517448501_1080;
   wire v3_1517448501_1081;
   wire v3_1517448501_1082;
   wire v3_1517448501_1083;
   wire v3_1517448501_1084;
   wire v3_1517448501_1085;
   wire v3_1517448501_1086;
   wire v3_1517448501_1087;
   wire v3_1517448501_1088;
   wire v3_1517448501_1089;
   wire v3_1517448501_1090;
   wire v3_1517448501_1091;
   wire v3_1517448501_1092;
   wire v3_1517448501_1093;
   wire v3_1517448501_1094;
   wire v3_1517448501_1095;
   wire v3_1517448501_1096;
   wire v3_1517448501_1097;
   wire v3_1517448501_1098;
   wire v3_1517448501_1099;
   wire v3_1517448501_1100;
   wire v3_1517448501_1101;
   wire v3_1517448501_1102;
   wire v3_1517448501_1103;
   wire v3_1517448501_1104;
   wire v3_1517448501_1105;
   wire v3_1517448501_1106;
   wire v3_1517448501_1107;
   wire v3_1517448501_1108;
   wire v3_1517448501_1109;
   wire v3_1517448501_1110;
   wire v3_1517448501_1111;
   wire v3_1517448501_1112;
   wire v3_1517448501_1113;
   wire v3_1517448501_1114;
   wire v3_1517448501_1115;
   wire v3_1517448501_1116;
   wire v3_1517448501_1117;
   wire v3_1517448501_1118;
   wire v3_1517448501_1119;
   wire v3_1517448501_1120;
   wire v3_1517448501_1121;
   wire v3_1517448501_1122;
   wire v3_1517448501_1123;
   wire v3_1517448501_1124;
   wire v3_1517448501_1125;
   wire v3_1517448501_1126;
   wire v3_1517448501_1127;
   wire v3_1517448501_1128;
   wire v3_1517448501_1129;
   wire v3_1517448501_1130;
   wire v3_1517448501_1131;
   wire v3_1517448501_1132;
   wire v3_1517448501_1133;
   wire v3_1517448501_1134;
   wire v3_1517448501_1135;
   wire v3_1517448501_1136;
   wire v3_1517448501_1137;
   wire v3_1517448501_1138;
   wire v3_1517448501_1139;
   wire v3_1517448501_1140;
   wire v3_1517448501_1141;
   wire v3_1517448501_1142;
   wire v3_1517448501_1143;
   wire v3_1517448501_1144;
   wire v3_1517448501_1145;
   wire v3_1517448501_1146;
   wire v3_1517448501_1147;
   wire v3_1517448501_1148;
   wire v3_1517448501_1149;
   wire v3_1517448501_1150;
   wire v3_1517448501_1151;
   wire v3_1517448501_1152;
   wire v3_1517448501_1153;
   wire v3_1517448501_1154;
   wire v3_1517448501_1155;
   wire v3_1517448501_1156;
   wire v3_1517448501_1157;
   wire v3_1517448501_1158;
   wire v3_1517448501_1159;
   wire v3_1517448501_1160;
   wire v3_1517448501_1161;
   wire v3_1517448501_1162;
   wire v3_1517448501_1163;
   wire v3_1517448501_1164;
   wire v3_1517448501_1165;
   wire v3_1517448501_1166;
   wire v3_1517448501_1167;
   wire v3_1517448501_1168;
   wire v3_1517448501_1169;
   wire v3_1517448501_1170;
   wire v3_1517448501_1171;
   wire v3_1517448501_1172;
   wire v3_1517448501_1173;
   wire v3_1517448501_1174;
   wire v3_1517448501_1175;
   wire v3_1517448501_1176;
   wire v3_1517448501_1177;
   wire v3_1517448501_1178;
   wire v3_1517448501_1179;
   wire v3_1517448501_1180;
   wire v3_1517448501_1181;
   wire v3_1517448501_1182;
   wire v3_1517448501_1183;
   wire v3_1517448501_1184;
   wire v3_1517448501_1185;
   wire v3_1517448501_1186;
   wire v3_1517448501_1187;
   wire v3_1517448501_1188;
   wire v3_1517448501_1189;
   wire v3_1517448501_1190;
   wire v3_1517448501_1191;
   wire v3_1517448501_1192;
   wire v3_1517448501_1193;
   wire v3_1517448501_1194;
   wire v3_1517448501_1195;
   wire v3_1517448501_1196;
   wire v3_1517448501_1197;
   wire v3_1517448501_1198;
   wire v3_1517448501_1199;
   wire v3_1517448501_1200;
   wire v3_1517448501_1201;
   wire v3_1517448501_1202;
   wire v3_1517448501_1203;
   wire v3_1517448501_1204;
   wire v3_1517448501_1205;
   wire v3_1517448501_1206;
   wire v3_1517448501_1207;
   wire v3_1517448501_1208;
   wire v3_1517448501_1209;
   wire v3_1517448501_1210;
   wire v3_1517448501_1211;
   wire v3_1517448501_1212;
   wire v3_1517448501_1213;
   wire v3_1517448501_1214;
   wire v3_1517448501_1215;
   wire v3_1517448501_1216;
   wire v3_1517448501_1217;
   wire v3_1517448501_1218;
   wire v3_1517448501_1219;
   wire v3_1517448501_1220;
   wire v3_1517448501_1221;
   wire v3_1517448501_1222;
   wire v3_1517448501_1223;
   wire v3_1517448501_1224;
   wire v3_1517448501_1225;
   wire v3_1517448501_1226;
   wire v3_1517448501_1227;
   wire v3_1517448501_1228;
   wire [7:0] v3_1517448501_1229;
   wire v3_1517448501_1230;
   wire v3_1517448501_1231;
   wire v3_1517448501_1232;
   wire v3_1517448501_1233;
   wire v3_1517448501_1234;
   wire v3_1517448501_1235;
   wire v3_1517448501_1236;
   wire v3_1517448501_1237;
   wire v3_1517448501_1238;
   wire v3_1517448501_1239;
   wire v3_1517448501_1240;
   wire v3_1517448501_1241;
   wire v3_1517448501_1242;
   wire v3_1517448501_1243;
   wire v3_1517448501_1244;
   wire v3_1517448501_1245;
   wire v3_1517448501_1246;
   wire v3_1517448501_1247;
   wire v3_1517448501_1248;
   wire v3_1517448501_1249;
   wire v3_1517448501_1250;
   wire v3_1517448501_1251;
   wire v3_1517448501_1252;
   wire v3_1517448501_1253;
   wire v3_1517448501_1254;
   wire v3_1517448501_1255;
   wire v3_1517448501_1256;
   wire v3_1517448501_1257;
   wire v3_1517448501_1258;
   wire v3_1517448501_1259;
   wire v3_1517448501_1260;
   wire v3_1517448501_1261;
   wire v3_1517448501_1262;
   wire v3_1517448501_1263;
   wire v3_1517448501_1264;
   wire v3_1517448501_1265;
   wire v3_1517448501_1266;
   wire v3_1517448501_1267;
   wire v3_1517448501_1268;
   wire v3_1517448501_1269;
   wire v3_1517448501_1270;
   wire v3_1517448501_1271;
   wire v3_1517448501_1272;
   wire v3_1517448501_1273;
   wire v3_1517448501_1274;
   wire v3_1517448501_1275;
   wire v3_1517448501_1276;
   wire v3_1517448501_1277;
   wire v3_1517448501_1278;
   wire v3_1517448501_1279;
   wire v3_1517448501_1280;
   wire v3_1517448501_1281;
   wire v3_1517448501_1282;
   wire v3_1517448501_1283;
   wire v3_1517448501_1284;
   wire v3_1517448501_1285;
   wire v3_1517448501_1286;
   wire v3_1517448501_1287;
   wire v3_1517448501_1288;
   wire v3_1517448501_1289;
   wire v3_1517448501_1290;
   wire v3_1517448501_1291;
   wire v3_1517448501_1292;
   wire v3_1517448501_1293;
   wire v3_1517448501_1294;
   wire v3_1517448501_1295;
   wire v3_1517448501_1296;
   wire v3_1517448501_1297;
   wire v3_1517448501_1298;
   wire v3_1517448501_1299;
   wire v3_1517448501_1300;
   wire v3_1517448501_1301;
   wire v3_1517448501_1302;
   wire v3_1517448501_1303;
   wire v3_1517448501_1304;
   wire v3_1517448501_1305;
   wire v3_1517448501_1306;
   wire v3_1517448501_1307;
   wire v3_1517448501_1308;
   wire v3_1517448501_1309;
   wire v3_1517448501_1310;
   wire v3_1517448501_1311;
   wire v3_1517448501_1312;
   wire v3_1517448501_1313;
   wire v3_1517448501_1314;
   wire v3_1517448501_1315;
   wire v3_1517448501_1316;
   wire v3_1517448501_1317;
   wire v3_1517448501_1318;
   wire v3_1517448501_1319;
   wire v3_1517448501_1320;
   wire v3_1517448501_1321;
   wire v3_1517448501_1322;
   wire v3_1517448501_1323;
   wire v3_1517448501_1324;
   wire v3_1517448501_1325;
   wire v3_1517448501_1326;
   wire v3_1517448501_1327;
   wire v3_1517448501_1328;
   wire v3_1517448501_1329;
   wire v3_1517448501_1330;
   wire v3_1517448501_1331;
   wire v3_1517448501_1332;
   wire v3_1517448501_1333;
   wire v3_1517448501_1334;
   wire v3_1517448501_1335;
   wire v3_1517448501_1336;
   wire v3_1517448501_1337;
   wire v3_1517448501_1338;
   wire v3_1517448501_1339;
   wire v3_1517448501_1340;
   wire v3_1517448501_1341;
   wire v3_1517448501_1342;
   wire v3_1517448501_1343;
   wire v3_1517448501_1344;
   wire v3_1517448501_1345;
   wire v3_1517448501_1346;
   wire v3_1517448501_1347;
   wire v3_1517448501_1348;
   wire v3_1517448501_1349;
   wire v3_1517448501_1350;
   wire v3_1517448501_1351;
   wire v3_1517448501_1352;
   wire v3_1517448501_1353;
   wire v3_1517448501_1354;
   wire v3_1517448501_1355;
   wire v3_1517448501_1356;
   wire v3_1517448501_1357;
   wire v3_1517448501_1358;
   wire v3_1517448501_1359;
   wire v3_1517448501_1360;
   wire v3_1517448501_1361;
   wire v3_1517448501_1362;
   wire v3_1517448501_1363;
   wire v3_1517448501_1364;
   wire v3_1517448501_1365;
   wire v3_1517448501_1366;
   wire v3_1517448501_1367;
   wire v3_1517448501_1368;
   wire v3_1517448501_1369;
   wire v3_1517448501_1370;
   wire v3_1517448501_1371;
   wire v3_1517448501_1372;
   wire v3_1517448501_1373;
   wire v3_1517448501_1374;
   wire v3_1517448501_1375;
   wire v3_1517448501_1376;
   wire v3_1517448501_1377;
   wire v3_1517448501_1378;
   wire v3_1517448501_1379;
   wire v3_1517448501_1380;
   wire v3_1517448501_1381;
   wire v3_1517448501_1382;
   wire v3_1517448501_1383;
   wire v3_1517448501_1384;
   wire v3_1517448501_1385;
   wire v3_1517448501_1386;
   wire v3_1517448501_1387;
   wire v3_1517448501_1388;
   wire v3_1517448501_1389;
   wire v3_1517448501_1390;
   wire v3_1517448501_1391;
   wire v3_1517448501_1392;
   wire v3_1517448501_1393;
   wire v3_1517448501_1394;
   wire v3_1517448501_1395;
   wire v3_1517448501_1396;
   wire v3_1517448501_1397;
   wire v3_1517448501_1398;
   wire v3_1517448501_1399;
   wire v3_1517448501_1400;
   wire v3_1517448501_1401;
   wire v3_1517448501_1402;
   wire v3_1517448501_1403;
   wire v3_1517448501_1404;
   wire v3_1517448501_1405;
   wire v3_1517448501_1406;
   wire v3_1517448501_1407;
   wire v3_1517448501_1408;
   wire v3_1517448501_1409;
   wire v3_1517448501_1410;
   wire v3_1517448501_1411;
   wire v3_1517448501_1412;
   wire v3_1517448501_1413;
   wire v3_1517448501_1414;
   wire v3_1517448501_1415;
   wire v3_1517448501_1416;
   wire v3_1517448501_1417;
   wire v3_1517448501_1418;
   wire v3_1517448501_1419;
   wire v3_1517448501_1420;
   wire v3_1517448501_1421;
   wire v3_1517448501_1422;
   wire v3_1517448501_1423;
   wire v3_1517448501_1424;
   wire v3_1517448501_1425;
   wire v3_1517448501_1426;
   wire v3_1517448501_1427;
   wire v3_1517448501_1428;
   wire v3_1517448501_1429;
   wire v3_1517448501_1430;
   wire v3_1517448501_1431;
   wire v3_1517448501_1432;
   wire v3_1517448501_1433;
   wire v3_1517448501_1434;
   wire v3_1517448501_1435;
   wire v3_1517448501_1436;
   wire v3_1517448501_1437;
   wire v3_1517448501_1438;
   wire v3_1517448501_1439;
   wire v3_1517448501_1440;
   wire v3_1517448501_1441;
   wire v3_1517448501_1442;
   wire v3_1517448501_1443;
   wire v3_1517448501_1444;
   wire v3_1517448501_1445;
   wire v3_1517448501_1446;
   wire v3_1517448501_1447;
   wire v3_1517448501_1448;
   wire v3_1517448501_1449;
   wire v3_1517448501_1450;
   wire v3_1517448501_1451;
   wire v3_1517448501_1452;
   wire v3_1517448501_1453;
   wire v3_1517448501_1454;
   wire v3_1517448501_1455;
   wire v3_1517448501_1456;
   wire v3_1517448501_1457;
   wire v3_1517448501_1458;
   wire v3_1517448501_1459;
   wire v3_1517448501_1460;
   wire v3_1517448501_1461;
   wire v3_1517448501_1462;
   wire v3_1517448501_1463;
   wire v3_1517448501_1464;
   wire v3_1517448501_1465;
   wire v3_1517448501_1466;
   wire v3_1517448501_1467;
   wire v3_1517448501_1468;
   wire v3_1517448501_1469;
   wire v3_1517448501_1470;
   wire v3_1517448501_1471;
   wire v3_1517448501_1472;
   wire v3_1517448501_1473;
   wire v3_1517448501_1474;
   wire v3_1517448501_1475;
   wire v3_1517448501_1476;
   wire v3_1517448501_1477;
   wire v3_1517448501_1478;
   wire v3_1517448501_1479;
   wire v3_1517448501_1480;
   wire v3_1517448501_1481;
   wire v3_1517448501_1482;
   wire v3_1517448501_1483;
   wire v3_1517448501_1484;
   wire v3_1517448501_1485;
   wire v3_1517448501_1486;
   wire v3_1517448501_1487;
   wire v3_1517448501_1488;
   wire v3_1517448501_1489;
   wire v3_1517448501_1490;
   wire v3_1517448501_1491;
   wire v3_1517448501_1492;
   wire v3_1517448501_1493;
   wire v3_1517448501_1494;
   wire v3_1517448501_1495;
   wire v3_1517448501_1496;
   wire v3_1517448501_1497;
   wire v3_1517448501_1498;
   wire v3_1517448501_1499;
   wire v3_1517448501_1500;
   wire v3_1517448501_1501;
   wire v3_1517448501_1502;
   wire v3_1517448501_1503;
   wire v3_1517448501_1504;
   wire v3_1517448501_1505;
   wire v3_1517448501_1506;
   wire v3_1517448501_1507;
   wire v3_1517448501_1508;
   wire v3_1517448501_1509;
   wire v3_1517448501_1510;
   wire v3_1517448501_1511;
   wire v3_1517448501_1512;
   wire v3_1517448501_1513;
   wire v3_1517448501_1514;
   wire v3_1517448501_1515;
   wire v3_1517448501_1516;
   wire v3_1517448501_1517;
   wire v3_1517448501_1518;
   wire v3_1517448501_1519;
   wire v3_1517448501_1520;
   wire v3_1517448501_1521;
   wire v3_1517448501_1522;
   wire v3_1517448501_1523;
   wire v3_1517448501_1524;
   wire v3_1517448501_1525;
   wire v3_1517448501_1526;
   wire v3_1517448501_1527;
   wire v3_1517448501_1528;
   wire v3_1517448501_1529;
   wire v3_1517448501_1530;
   wire v3_1517448501_1531;
   wire v3_1517448501_1532;
   wire v3_1517448501_1533;
   wire v3_1517448501_1534;
   wire v3_1517448501_1535;
   wire v3_1517448501_1536;
   wire v3_1517448501_1537;
   wire v3_1517448501_1538;
   wire v3_1517448501_1539;
   wire v3_1517448501_1540;
   wire v3_1517448501_1541;
   wire v3_1517448501_1542;
   wire v3_1517448501_1543;
   wire v3_1517448501_1544;
   wire v3_1517448501_1545;
   wire v3_1517448501_1546;
   wire v3_1517448501_1547;
   wire v3_1517448501_1548;
   wire v3_1517448501_1549;
   wire v3_1517448501_1550;
   wire v3_1517448501_1551;
   wire v3_1517448501_1552;
   wire v3_1517448501_1553;
   wire v3_1517448501_1554;
   wire v3_1517448501_1555;
   wire v3_1517448501_1556;
   wire v3_1517448501_1557;
   wire v3_1517448501_1558;
   wire v3_1517448501_1559;
   wire v3_1517448501_1560;
   wire v3_1517448501_1561;
   wire v3_1517448501_1562;
   wire v3_1517448501_1563;
   wire v3_1517448501_1564;
   wire v3_1517448501_1565;
   wire v3_1517448501_1566;
   wire v3_1517448501_1567;
   wire v3_1517448501_1568;
   wire v3_1517448501_1569;
   wire v3_1517448501_1570;
   wire v3_1517448501_1571;
   wire v3_1517448501_1572;
   wire v3_1517448501_1573;
   wire v3_1517448501_1574;
   wire v3_1517448501_1575;
   wire v3_1517448501_1576;
   wire v3_1517448501_1577;
   wire v3_1517448501_1578;
   wire v3_1517448501_1579;
   wire v3_1517448501_1580;
   wire v3_1517448501_1581;
   wire v3_1517448501_1582;
   wire v3_1517448501_1583;
   wire v3_1517448501_1584;
   wire v3_1517448501_1585;
   wire v3_1517448501_1586;
   wire v3_1517448501_1587;
   wire v3_1517448501_1588;
   wire v3_1517448501_1589;
   wire v3_1517448501_1590;
   wire v3_1517448501_1591;
   wire v3_1517448501_1592;
   wire v3_1517448501_1593;
   wire v3_1517448501_1594;
   wire v3_1517448501_1595;
   wire v3_1517448501_1596;
   wire v3_1517448501_1597;
   wire v3_1517448501_1598;
   wire v3_1517448501_1599;
   wire v3_1517448501_1600;
   wire v3_1517448501_1601;
   wire v3_1517448501_1602;
   wire v3_1517448501_1603;
   wire v3_1517448501_1604;
   wire v3_1517448501_1605;
   wire v3_1517448501_1606;
   wire v3_1517448501_1607;
   wire v3_1517448501_1608;
   wire v3_1517448501_1609;
   wire v3_1517448501_1610;
   wire v3_1517448501_1611;
   wire v3_1517448501_1612;
   wire v3_1517448501_1613;
   wire v3_1517448501_1614;
   wire v3_1517448501_1615;
   wire v3_1517448501_1616;
   wire v3_1517448501_1617;
   wire v3_1517448501_1618;
   wire v3_1517448501_1619;
   wire v3_1517448501_1620;
   wire v3_1517448501_1621;
   wire v3_1517448501_1622;
   wire v3_1517448501_1623;
   wire v3_1517448501_1624;
   wire v3_1517448501_1625;
   wire v3_1517448501_1626;
   wire v3_1517448501_1627;
   wire v3_1517448501_1628;
   wire v3_1517448501_1629;
   wire v3_1517448501_1630;
   wire v3_1517448501_1631;
   wire v3_1517448501_1632;
   wire v3_1517448501_1633;
   wire v3_1517448501_1634;
   wire v3_1517448501_1635;
   wire v3_1517448501_1636;
   wire v3_1517448501_1637;
   wire v3_1517448501_1638;
   wire v3_1517448501_1639;
   wire v3_1517448501_1640;
   wire v3_1517448501_1641;
   wire v3_1517448501_1642;
   wire v3_1517448501_1643;
   wire v3_1517448501_1644;
   wire v3_1517448501_1645;
   wire v3_1517448501_1646;
   wire v3_1517448501_1647;
   wire v3_1517448501_1648;
   wire v3_1517448501_1649;
   wire v3_1517448501_1650;
   wire v3_1517448501_1651;
   wire v3_1517448501_1652;
   wire v3_1517448501_1653;
   wire v3_1517448501_1654;
   wire v3_1517448501_1655;
   wire v3_1517448501_1656;
   wire v3_1517448501_1657;
   wire v3_1517448501_1658;
   wire v3_1517448501_1659;
   wire v3_1517448501_1660;
   wire v3_1517448501_1661;
   wire v3_1517448501_1662;
   wire v3_1517448501_1663;
   wire v3_1517448501_1664;
   wire v3_1517448501_1665;
   wire v3_1517448501_1666;
   wire v3_1517448501_1667;
   wire v3_1517448501_1668;
   wire v3_1517448501_1669;
   wire v3_1517448501_1670;
   wire v3_1517448501_1671;
   wire v3_1517448501_1672;
   wire v3_1517448501_1673;
   wire v3_1517448501_1674;
   wire v3_1517448501_1675;
   wire v3_1517448501_1676;
   wire v3_1517448501_1677;
   wire v3_1517448501_1678;
   wire v3_1517448501_1679;
   wire v3_1517448501_1680;
   wire v3_1517448501_1681;
   wire v3_1517448501_1682;
   wire v3_1517448501_1683;
   wire v3_1517448501_1684;
   wire v3_1517448501_1685;
   wire v3_1517448501_1686;
   wire v3_1517448501_1687;
   wire v3_1517448501_1688;
   wire v3_1517448501_1689;
   wire v3_1517448501_1690;
   wire v3_1517448501_1691;
   wire v3_1517448501_1692;
   wire v3_1517448501_1693;
   wire v3_1517448501_1694;
   wire v3_1517448501_1695;
   wire v3_1517448501_1696;
   wire v3_1517448501_1697;
   wire v3_1517448501_1698;
   wire v3_1517448501_1699;
   wire v3_1517448501_1700;
   wire v3_1517448501_1701;
   wire v3_1517448501_1702;
   wire v3_1517448501_1703;
   wire v3_1517448501_1704;
   wire v3_1517448501_1705;
   wire v3_1517448501_1706;
   wire v3_1517448501_1707;
   wire v3_1517448501_1708;
   wire v3_1517448501_1709;
   wire v3_1517448501_1710;
   wire v3_1517448501_1711;
   wire v3_1517448501_1712;
   wire v3_1517448501_1713;
   wire v3_1517448501_1714;
   wire v3_1517448501_1715;
   wire v3_1517448501_1716;
   wire v3_1517448501_1717;
   wire v3_1517448501_1718;
   wire v3_1517448501_1719;
   wire v3_1517448501_1720;
   wire v3_1517448501_1721;
   wire v3_1517448501_1722;
   wire v3_1517448501_1723;
   wire v3_1517448501_1724;
   wire v3_1517448501_1725;
   wire v3_1517448501_1726;
   wire v3_1517448501_1727;
   wire v3_1517448501_1728;
   wire v3_1517448501_1729;
   wire v3_1517448501_1730;
   wire v3_1517448501_1731;
   wire v3_1517448501_1732;
   wire v3_1517448501_1733;
   wire v3_1517448501_1734;
   wire v3_1517448501_1735;
   wire v3_1517448501_1736;
   wire v3_1517448501_1737;
   wire v3_1517448501_1738;
   wire v3_1517448501_1739;
   wire v3_1517448501_1740;
   wire v3_1517448501_1741;
   wire v3_1517448501_1742;
   wire v3_1517448501_1743;
   wire v3_1517448501_1744;
   wire v3_1517448501_1745;
   wire v3_1517448501_1746;
   wire v3_1517448501_1747;
   wire v3_1517448501_1748;
   wire v3_1517448501_1749;
   wire v3_1517448501_1750;
   wire v3_1517448501_1751;
   wire v3_1517448501_1752;
   wire v3_1517448501_1753;
   wire v3_1517448501_1754;
   wire v3_1517448501_1755;
   wire v3_1517448501_1756;
   wire v3_1517448501_1757;
   wire v3_1517448501_1758;
   wire v3_1517448501_1759;
   wire v3_1517448501_1760;
   wire v3_1517448501_1761;
   wire v3_1517448501_1762;
   wire v3_1517448501_1763;
   wire v3_1517448501_1764;
   wire v3_1517448501_1765;
   wire v3_1517448501_1766;
   wire v3_1517448501_1767;
   wire v3_1517448501_1768;
   wire v3_1517448501_1769;
   wire v3_1517448501_1770;
   wire v3_1517448501_1771;
   wire v3_1517448501_1772;
   wire v3_1517448501_1773;
   wire v3_1517448501_1774;
   wire v3_1517448501_1775;
   wire v3_1517448501_1776;
   wire v3_1517448501_1777;
   wire v3_1517448501_1778;
   wire v3_1517448501_1779;
   wire v3_1517448501_1780;
   wire v3_1517448501_1781;
   wire v3_1517448501_1782;
   wire v3_1517448501_1783;
   wire v3_1517448501_1784;
   wire v3_1517448501_1785;
   wire v3_1517448501_1786;
   wire v3_1517448501_1787;
   wire v3_1517448501_1788;
   wire v3_1517448501_1789;
   wire v3_1517448501_1790;
   wire v3_1517448501_1791;
   wire v3_1517448501_1792;
   wire v3_1517448501_1793;
   wire v3_1517448501_1794;
   wire v3_1517448501_1795;
   wire v3_1517448501_1796;
   wire v3_1517448501_1797;
   wire v3_1517448501_1798;
   wire v3_1517448501_1799;
   wire v3_1517448501_1800;
   wire v3_1517448501_1801;
   wire v3_1517448501_1802;
   wire v3_1517448501_1803;
   wire v3_1517448501_1804;
   wire v3_1517448501_1805;
   wire v3_1517448501_1806;
   wire v3_1517448501_1807;
   wire v3_1517448501_1808;
   wire v3_1517448501_1809;
   wire v3_1517448501_1810;
   wire v3_1517448501_1811;
   wire v3_1517448501_1812;
   wire v3_1517448501_1813;
   wire v3_1517448501_1814;
   wire v3_1517448501_1815;
   wire v3_1517448501_1816;
   wire v3_1517448501_1817;
   wire v3_1517448501_1818;
   wire v3_1517448501_1819;
   wire v3_1517448501_1820;
   wire v3_1517448501_1821;
   wire v3_1517448501_1822;
   wire v3_1517448501_1823;
   wire v3_1517448501_1824;
   wire v3_1517448501_1825;
   wire v3_1517448501_1826;
   wire v3_1517448501_1827;
   wire v3_1517448501_1828;
   wire v3_1517448501_1829;
   wire v3_1517448501_1830;
   wire v3_1517448501_1831;
   wire v3_1517448501_1832;
   wire v3_1517448501_1833;
   wire v3_1517448501_1834;
   wire v3_1517448501_1835;
   wire v3_1517448501_1836;
   wire v3_1517448501_1837;
   wire v3_1517448501_1838;
   wire v3_1517448501_1839;
   wire v3_1517448501_1840;
   wire v3_1517448501_1841;
   wire v3_1517448501_1842;
   wire v3_1517448501_1843;
   wire v3_1517448501_1844;
   wire v3_1517448501_1845;
   wire v3_1517448501_1846;
   wire v3_1517448501_1847;
   wire v3_1517448501_1848;
   wire v3_1517448501_1849;
   wire v3_1517448501_1850;
   wire v3_1517448501_1851;
   wire v3_1517448501_1852;
   wire v3_1517448501_1853;
   wire v3_1517448501_1854;
   wire v3_1517448501_1855;
   wire v3_1517448501_1856;
   wire v3_1517448501_1857;
   wire v3_1517448501_1858;
   wire v3_1517448501_1859;
   wire v3_1517448501_1860;
   wire v3_1517448501_1861;
   wire v3_1517448501_1862;
   wire v3_1517448501_1863;
   wire v3_1517448501_1864;
   wire v3_1517448501_1865;
   wire v3_1517448501_1866;
   wire v3_1517448501_1867;
   wire v3_1517448501_1868;
   wire v3_1517448501_1869;
   wire v3_1517448501_1870;
   wire v3_1517448501_1871;
   wire v3_1517448501_1872;
   wire v3_1517448501_1873;
   wire v3_1517448501_1874;
   wire v3_1517448501_1875;
   wire v3_1517448501_1876;
   wire v3_1517448501_1877;
   wire v3_1517448501_1878;
   wire v3_1517448501_1879;
   wire v3_1517448501_1880;
   wire v3_1517448501_1881;
   wire v3_1517448501_1882;
   wire v3_1517448501_1883;
   wire v3_1517448501_1884;
   wire v3_1517448501_1885;
   wire v3_1517448501_1886;
   wire v3_1517448501_1887;
   wire v3_1517448501_1888;
   wire v3_1517448501_1889;
   wire v3_1517448501_1890;
   wire v3_1517448501_1891;
   wire v3_1517448501_1892;
   wire v3_1517448501_1893;
   wire v3_1517448501_1894;
   wire v3_1517448501_1895;
   wire v3_1517448501_1896;
   wire v3_1517448501_1897;
   wire v3_1517448501_1898;
   wire v3_1517448501_1899;
   wire v3_1517448501_1900;
   wire v3_1517448501_1901;
   wire v3_1517448501_1902;
   wire v3_1517448501_1903;
   wire v3_1517448501_1904;
   wire v3_1517448501_1905;
   wire v3_1517448501_1906;
   wire v3_1517448501_1907;
   wire v3_1517448501_1908;
   wire v3_1517448501_1909;
   wire v3_1517448501_1910;
   wire v3_1517448501_1911;
   wire v3_1517448501_1912;
   wire v3_1517448501_1913;
   wire v3_1517448501_1914;
   wire v3_1517448501_1915;
   wire v3_1517448501_1916;
   wire v3_1517448501_1917;
   wire v3_1517448501_1918;
   wire v3_1517448501_1919;
   wire v3_1517448501_1920;
   wire v3_1517448501_1921;
   wire v3_1517448501_1922;
   wire v3_1517448501_1923;
   wire v3_1517448501_1924;
   wire v3_1517448501_1925;
   wire v3_1517448501_1926;
   wire v3_1517448501_1927;
   wire v3_1517448501_1928;
   wire v3_1517448501_1929;
   wire v3_1517448501_1930;
   wire v3_1517448501_1931;
   wire v3_1517448501_1932;
   wire v3_1517448501_1933;
   wire v3_1517448501_1934;
   wire v3_1517448501_1935;
   wire v3_1517448501_1936;
   wire v3_1517448501_1937;
   wire v3_1517448501_1938;
   wire v3_1517448501_1939;
   wire v3_1517448501_1940;
   wire v3_1517448501_1941;
   wire v3_1517448501_1942;
   wire v3_1517448501_1943;
   wire v3_1517448501_1944;
   wire v3_1517448501_1945;
   wire v3_1517448501_1946;
   wire v3_1517448501_1947;
   wire v3_1517448501_1948;
   wire v3_1517448501_1949;
   wire v3_1517448501_1950;
   wire v3_1517448501_1951;
   wire v3_1517448501_1952;
   wire v3_1517448501_1953;
   wire v3_1517448501_1954;
   wire v3_1517448501_1955;
   wire v3_1517448501_1956;
   wire v3_1517448501_1957;
   wire v3_1517448501_1958;
   wire v3_1517448501_1959;
   wire v3_1517448501_1960;
   wire v3_1517448501_1961;
   wire v3_1517448501_1962;
   wire v3_1517448501_1963;
   wire v3_1517448501_1964;
   wire v3_1517448501_1965;
   wire v3_1517448501_1966;
   wire v3_1517448501_1967;
   wire v3_1517448501_1968;
   wire v3_1517448501_1969;
   wire v3_1517448501_1970;
   wire v3_1517448501_1971;
   wire v3_1517448501_1972;
   wire v3_1517448501_1973;
   wire v3_1517448501_1974;
   wire v3_1517448501_1975;
   wire v3_1517448501_1976;
   wire v3_1517448501_1977;
   wire v3_1517448501_1978;
   wire v3_1517448501_1979;
   wire v3_1517448501_1980;
   wire v3_1517448501_1981;
   wire v3_1517448501_1982;
   wire v3_1517448501_1983;
   wire v3_1517448501_1984;
   wire v3_1517448501_1985;
   wire v3_1517448501_1986;
   wire v3_1517448501_1987;
   wire v3_1517448501_1988;
   wire v3_1517448501_1989;
   wire v3_1517448501_1990;
   wire v3_1517448501_1991;
   wire v3_1517448501_1992;
   wire v3_1517448501_1993;
   wire v3_1517448501_1994;
   wire v3_1517448501_1995;
   wire v3_1517448501_1996;
   wire v3_1517448501_1997;
   wire v3_1517448501_1998;
   wire v3_1517448501_1999;
   wire v3_1517448501_2000;
   wire v3_1517448501_2001;
   wire v3_1517448501_2002;
   wire v3_1517448501_2003;
   wire v3_1517448501_2004;
   wire v3_1517448501_2005;
   wire v3_1517448501_2006;
   wire v3_1517448501_2007;
   wire v3_1517448501_2008;
   wire v3_1517448501_2009;
   wire v3_1517448501_2010;
   wire v3_1517448501_2011;
   wire v3_1517448501_2012;
   wire v3_1517448501_2013;
   wire v3_1517448501_2014;
   wire v3_1517448501_2015;
   wire v3_1517448501_2016;
   wire v3_1517448501_2017;
   wire v3_1517448501_2018;
   wire v3_1517448501_2019;
   wire v3_1517448501_2020;
   wire v3_1517448501_2021;
   wire v3_1517448501_2022;
   wire v3_1517448501_2023;
   wire v3_1517448501_2024;
   wire v3_1517448501_2025;
   wire v3_1517448501_2026;
   wire v3_1517448501_2027;
   wire v3_1517448501_2028;
   wire v3_1517448501_2029;
   wire v3_1517448501_2030;
   wire v3_1517448501_2031;
   wire v3_1517448501_2032;
   wire v3_1517448501_2033;
   wire v3_1517448501_2034;
   wire v3_1517448501_2035;
   wire v3_1517448501_2036;
   wire v3_1517448501_2037;
   wire v3_1517448501_2038;
   wire v3_1517448501_2039;
   wire v3_1517448501_2040;
   wire v3_1517448501_2041;
   wire v3_1517448501_2042;
   wire v3_1517448501_2043;
   wire v3_1517448501_2044;
   wire v3_1517448501_2045;
   wire v3_1517448501_2046;
   wire v3_1517448501_2047;
   wire v3_1517448501_2048;
   wire v3_1517448501_2049;
   wire v3_1517448501_2050;
   wire v3_1517448501_2051;
   wire v3_1517448501_2052;
   wire v3_1517448501_2053;
   wire v3_1517448501_2054;
   wire v3_1517448501_2055;
   wire v3_1517448501_2056;
   wire v3_1517448501_2057;
   wire v3_1517448501_2058;
   wire v3_1517448501_2059;
   wire v3_1517448501_2060;
   wire v3_1517448501_2061;
   wire v3_1517448501_2062;
   wire v3_1517448501_2063;
   wire v3_1517448501_2064;
   wire v3_1517448501_2065;
   wire v3_1517448501_2066;
   wire v3_1517448501_2067;
   wire v3_1517448501_2068;
   wire v3_1517448501_2069;
   wire v3_1517448501_2070;
   wire v3_1517448501_2071;
   wire v3_1517448501_2072;
   wire v3_1517448501_2073;
   wire v3_1517448501_2074;
   wire v3_1517448501_2075;
   wire v3_1517448501_2076;
   wire v3_1517448501_2077;
   wire v3_1517448501_2078;
   wire v3_1517448501_2079;
   wire v3_1517448501_2080;
   wire v3_1517448501_2081;
   wire v3_1517448501_2082;
   wire v3_1517448501_2083;
   wire v3_1517448501_2084;
   wire v3_1517448501_2085;
   wire v3_1517448501_2086;
   wire v3_1517448501_2087;
   wire v3_1517448501_2088;
   wire v3_1517448501_2089;
   wire v3_1517448501_2090;
   wire v3_1517448501_2091;
   wire v3_1517448501_2092;
   wire v3_1517448501_2093;
   wire v3_1517448501_2094;
   wire v3_1517448501_2095;
   wire v3_1517448501_2096;
   wire v3_1517448501_2097;
   wire v3_1517448501_2098;
   wire v3_1517448501_2099;
   wire v3_1517448501_2100;
   wire v3_1517448501_2101;
   wire v3_1517448501_2102;
   wire v3_1517448501_2103;
   wire v3_1517448501_2104;
   wire v3_1517448501_2105;
   wire v3_1517448501_2106;
   wire v3_1517448501_2107;
   wire v3_1517448501_2108;
   wire v3_1517448501_2109;
   wire v3_1517448501_2110;
   wire v3_1517448501_2111;
   wire v3_1517448501_2112;
   wire v3_1517448501_2113;
   wire v3_1517448501_2114;
   wire v3_1517448501_2115;
   wire v3_1517448501_2116;
   wire v3_1517448501_2117;
   wire v3_1517448501_2118;
   wire v3_1517448501_2119;
   wire v3_1517448501_2120;
   wire v3_1517448501_2121;
   wire v3_1517448501_2122;
   wire v3_1517448501_2123;
   wire v3_1517448501_2124;
   wire v3_1517448501_2125;
   wire v3_1517448501_2126;
   wire v3_1517448501_2127;
   wire v3_1517448501_2128;
   wire v3_1517448501_2129;
   wire v3_1517448501_2130;
   wire v3_1517448501_2131;
   wire v3_1517448501_2132;
   wire v3_1517448501_2133;
   wire v3_1517448501_2134;
   wire v3_1517448501_2135;
   wire v3_1517448501_2136;
   wire v3_1517448501_2137;
   wire v3_1517448501_2138;
   wire v3_1517448501_2139;
   wire v3_1517448501_2140;
   wire v3_1517448501_2141;
   wire v3_1517448501_2142;
   wire v3_1517448501_2143;
   wire v3_1517448501_2144;

   // Output Net Declarations
   wire id60;

   // Combinational Assignments
   assign id0 = 1'b0; 
   assign v3_1517448501_52 = 32'b00000000_00000000_00000000_00000111; 
   assign v3_1517448501_53 = 16'b00000000_00000000; 
   assign v3_1517448501_54 = {v_party_responder_0, v3_1517448501_53};
   assign v3_1517448501_55 = 5'b10000; 
   assign v3_1517448501_56 = v3_1517448501_59 ? ~v3_1517448501_58 : v3_1517448501_57;
   assign v3_1517448501_57 = v3_1517448501_54 >> v3_1517448501_55;
   assign v3_1517448501_58 = ~v3_1517448501_54 >> v3_1517448501_55;
   assign v3_1517448501_59 = v3_1517448501_54[31];
   assign v3_1517448501_60 = v3_1517448501_52 == v3_1517448501_56;
   assign v3_1517448501_61 = a_finished_responder_0 & v3_1517448501_60;
   assign v3_1517448501_62 = ~dve_invalid & v3_1517448501_61;
   assign v3_1517448501_64 = 16'b00000110_11101011; 
   assign v3_1517448501_66 = 16'b00000110_01100100; 
   assign v3_1517448501_68 = 16'b00000110_00110111; 
   assign v3_1517448501_70 = 32'b00000000_00000000_00000000_01001011; 
   assign v3_1517448501_71 = {v_party_nonce_responder_1, v3_1517448501_53};
   assign v3_1517448501_72 = v3_1517448501_75 ? ~v3_1517448501_74 : v3_1517448501_73;
   assign v3_1517448501_73 = v3_1517448501_71 >> v3_1517448501_55;
   assign v3_1517448501_74 = ~v3_1517448501_71 >> v3_1517448501_55;
   assign v3_1517448501_75 = v3_1517448501_71[31];
   assign v3_1517448501_76 = v3_1517448501_70 + v3_1517448501_72;
   assign v3_1517448501_77 = 32'b00000000_00000000_00000000_00001111; 
   assign v3_1517448501_78 = {v_party_responder_1, v3_1517448501_53};
   assign v3_1517448501_79 = v3_1517448501_82 ? ~v3_1517448501_81 : v3_1517448501_80;
   assign v3_1517448501_80 = v3_1517448501_78 >> v3_1517448501_55;
   assign v3_1517448501_81 = ~v3_1517448501_78 >> v3_1517448501_55;
   assign v3_1517448501_82 = v3_1517448501_78[31];
   assign v3_1517448501_83 = v3_1517448501_77 * v3_1517448501_79;
   assign v3_1517448501_84 = v3_1517448501_77 * v3_1517448501_83;
   assign v3_1517448501_85 = v3_1517448501_76 + v3_1517448501_84;
   assign v3_1517448501_86 = v3_1517448501_85[15:0];
   assign v3_1517448501_88 = 32'b00000000_00000000_00000000_00111100; 
   assign v3_1517448501_89 = {v_party_nonce_responder_0, v3_1517448501_53};
   assign v3_1517448501_90 = v3_1517448501_93 ? ~v3_1517448501_92 : v3_1517448501_91;
   assign v3_1517448501_91 = v3_1517448501_89 >> v3_1517448501_55;
   assign v3_1517448501_92 = ~v3_1517448501_89 >> v3_1517448501_55;
   assign v3_1517448501_93 = v3_1517448501_89[31];
   assign v3_1517448501_94 = v3_1517448501_88 + v3_1517448501_90;
   assign v3_1517448501_95 = v3_1517448501_77 * v3_1517448501_56;
   assign v3_1517448501_96 = v3_1517448501_77 * v3_1517448501_95;
   assign v3_1517448501_97 = v3_1517448501_94 + v3_1517448501_96;
   assign v3_1517448501_98 = v3_1517448501_97[15:0];
   assign v3_1517448501_99 = f78 ? v3_1517448501_98 : v_m_initiator_0;
   assign v3_1517448501_100 = f81 ? v3_1517448501_86 : v3_1517448501_99;
   assign v3_1517448501_101 = f84 ? v3_1517448501_68 : v3_1517448501_100;
   assign v3_1517448501_102 = f86 ? v3_1517448501_66 : v3_1517448501_101;
   assign v3_1517448501_103 = f88 ? v3_1517448501_64 : v3_1517448501_102;
   assign v3_1517448501_104 = 16'b00000000_00000000; 
   assign v3_1517448501_106 = {v_m_initiator_0, v3_1517448501_53};
   assign v3_1517448501_107 = v3_1517448501_110 ? ~v3_1517448501_109 : v3_1517448501_108;
   assign v3_1517448501_108 = v3_1517448501_106 >> v3_1517448501_55;
   assign v3_1517448501_109 = ~v3_1517448501_106 >> v3_1517448501_55;
   assign v3_1517448501_110 = v3_1517448501_106[31];
   assign v3_1517448501_111 = 32'b00000000_00000000_00000000_11100001; 
   assign v3_1517448501_112 = v3_1517448501_113 ? v3_1517448501_121 : v3_1517448501_120;
   assign v3_1517448501_113 = v3_1517448501_107[31];
   assign v3_1517448501_114 = v3_1517448501_111[31];
   assign v3_1517448501_115 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_116 = ~v3_1517448501_107 + v3_1517448501_115;
   assign v3_1517448501_117 = ~v3_1517448501_111 + v3_1517448501_115;
   assign v3_1517448501_118 = v3_1517448501_113 ? v3_1517448501_116 : v3_1517448501_107;
   assign v3_1517448501_119 = v3_1517448501_114 ? v3_1517448501_117 : v3_1517448501_111;
   assign v3_1517448501_120 = v3_1517448501_118 % v3_1517448501_119;
   assign v3_1517448501_121 = ~v3_1517448501_120 + v3_1517448501_115;
   assign v3_1517448501_122 = v3_1517448501_125 ? v3_1517448501_132 : v3_1517448501_131;
   assign v3_1517448501_123 = v3_1517448501_112[31];
   assign v3_1517448501_124 = v3_1517448501_77[31];
   assign v3_1517448501_125 = v3_1517448501_123 ^ v3_1517448501_124;
   assign v3_1517448501_126 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_127 = ~v3_1517448501_112 + v3_1517448501_126;
   assign v3_1517448501_128 = ~v3_1517448501_77 + v3_1517448501_126;
   assign v3_1517448501_129 = v3_1517448501_123 ? v3_1517448501_127 : v3_1517448501_112;
   assign v3_1517448501_130 = v3_1517448501_124 ? v3_1517448501_128 : v3_1517448501_77;
   assign v3_1517448501_131 = v3_1517448501_129 / v3_1517448501_130;
   assign v3_1517448501_132 = ~v3_1517448501_131 + v3_1517448501_126;
   assign v3_1517448501_133 = v3_1517448501_122[15:0];
   assign v3_1517448501_134 = f00 ? v3_1517448501_133 : v_party_nonce_initiator_0;
   assign v3_1517448501_135 = 16'b00000000_00000000; 
   assign v3_1517448501_141 = f79 ? v3_1517448501_98 : v_m_initiator_1;
   assign v3_1517448501_142 = f82 ? v3_1517448501_86 : v3_1517448501_141;
   assign v3_1517448501_143 = f85 ? v3_1517448501_68 : v3_1517448501_142;
   assign v3_1517448501_144 = f87 ? v3_1517448501_66 : v3_1517448501_143;
   assign v3_1517448501_145 = f89 ? v3_1517448501_64 : v3_1517448501_144;
   assign v3_1517448501_146 = 16'b00000000_00000000; 
   assign v3_1517448501_148 = {v_m_initiator_1, v3_1517448501_53};
   assign v3_1517448501_149 = v3_1517448501_152 ? ~v3_1517448501_151 : v3_1517448501_150;
   assign v3_1517448501_150 = v3_1517448501_148 >> v3_1517448501_55;
   assign v3_1517448501_151 = ~v3_1517448501_148 >> v3_1517448501_55;
   assign v3_1517448501_152 = v3_1517448501_148[31];
   assign v3_1517448501_153 = v3_1517448501_154 ? v3_1517448501_162 : v3_1517448501_161;
   assign v3_1517448501_154 = v3_1517448501_149[31];
   assign v3_1517448501_155 = v3_1517448501_111[31];
   assign v3_1517448501_156 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_157 = ~v3_1517448501_149 + v3_1517448501_156;
   assign v3_1517448501_158 = ~v3_1517448501_111 + v3_1517448501_156;
   assign v3_1517448501_159 = v3_1517448501_154 ? v3_1517448501_157 : v3_1517448501_149;
   assign v3_1517448501_160 = v3_1517448501_155 ? v3_1517448501_158 : v3_1517448501_111;
   assign v3_1517448501_161 = v3_1517448501_159 % v3_1517448501_160;
   assign v3_1517448501_162 = ~v3_1517448501_161 + v3_1517448501_156;
   assign v3_1517448501_163 = v3_1517448501_166 ? v3_1517448501_173 : v3_1517448501_172;
   assign v3_1517448501_164 = v3_1517448501_153[31];
   assign v3_1517448501_165 = v3_1517448501_77[31];
   assign v3_1517448501_166 = v3_1517448501_164 ^ v3_1517448501_165;
   assign v3_1517448501_167 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_168 = ~v3_1517448501_153 + v3_1517448501_167;
   assign v3_1517448501_169 = ~v3_1517448501_77 + v3_1517448501_167;
   assign v3_1517448501_170 = v3_1517448501_164 ? v3_1517448501_168 : v3_1517448501_153;
   assign v3_1517448501_171 = v3_1517448501_165 ? v3_1517448501_169 : v3_1517448501_77;
   assign v3_1517448501_172 = v3_1517448501_170 / v3_1517448501_171;
   assign v3_1517448501_173 = ~v3_1517448501_172 + v3_1517448501_167;
   assign v3_1517448501_174 = v3_1517448501_163[15:0];
   assign v3_1517448501_175 = f02 ? v3_1517448501_174 : v_party_nonce_initiator_1;
   assign v3_1517448501_176 = 16'b00000000_00000000; 
   assign v3_1517448501_178 = 16'b00000000_10011010; 
   assign v3_1517448501_180 = 32'b00000000_00000000_00000000_10100101; 
   assign v3_1517448501_181 = {v_party_nonce_initiator_1, v3_1517448501_53};
   assign v3_1517448501_182 = v3_1517448501_185 ? ~v3_1517448501_184 : v3_1517448501_183;
   assign v3_1517448501_183 = v3_1517448501_181 >> v3_1517448501_55;
   assign v3_1517448501_184 = ~v3_1517448501_181 >> v3_1517448501_55;
   assign v3_1517448501_185 = v3_1517448501_181[31];
   assign v3_1517448501_186 = v3_1517448501_180 + v3_1517448501_182;
   assign v3_1517448501_187 = v3_1517448501_186[15:0];
   assign v3_1517448501_189 = 32'b00000000_00000000_00000000_10010110; 
   assign v3_1517448501_190 = {v_party_nonce_initiator_0, v3_1517448501_53};
   assign v3_1517448501_191 = v3_1517448501_194 ? ~v3_1517448501_193 : v3_1517448501_192;
   assign v3_1517448501_192 = v3_1517448501_190 >> v3_1517448501_55;
   assign v3_1517448501_193 = ~v3_1517448501_190 >> v3_1517448501_55;
   assign v3_1517448501_194 = v3_1517448501_190[31];
   assign v3_1517448501_195 = v3_1517448501_189 + v3_1517448501_191;
   assign v3_1517448501_196 = v3_1517448501_195[15:0];
   assign v3_1517448501_198 = 16'b00001000_11101100; 
   assign v3_1517448501_200 = 16'b00001001_01100100; 
   assign v3_1517448501_202 = 16'b00001001_00110111; 
   assign v3_1517448501_204 = 16'b00001000_11101001; 
   assign v3_1517448501_206 = 16'b00001001_01100001; 
   assign v3_1517448501_208 = 16'b00001001_00110100; 
   assign v3_1517448501_210 = 16'b00000110_01000110; 
   assign v3_1517448501_212 = 16'b00000110_10111110; 
   assign v3_1517448501_214 = 16'b00000110_10010001; 
   assign v3_1517448501_216 = 16'b00001000_11101010; 
   assign v3_1517448501_218 = 16'b00001001_01100010; 
   assign v3_1517448501_220 = 16'b00001001_00110101; 
   assign v3_1517448501_222 = 16'b00001000_11110010; 
   assign v3_1517448501_224 = 16'b00001001_01101010; 
   assign v3_1517448501_226 = 16'b00001001_00111101; 
   assign v3_1517448501_228 = 16'b00001000_11101111; 
   assign v3_1517448501_230 = 16'b00001001_01100111; 
   assign v3_1517448501_232 = 16'b00001001_00111010; 
   assign v3_1517448501_234 = 16'b00001000_11110101; 
   assign v3_1517448501_236 = 16'b00001001_01101101; 
   assign v3_1517448501_238 = 16'b00001001_01000000; 
   assign v3_1517448501_240 = 16'b00001010_00100101; 
   assign v3_1517448501_242 = f30 ? v3_1517448501_208 : v_m_responder_0;
   assign v3_1517448501_243 = f33 ? v3_1517448501_240 : v3_1517448501_242;
   assign v3_1517448501_244 = f36 ? v3_1517448501_238 : v3_1517448501_243;
   assign v3_1517448501_245 = f38 ? v3_1517448501_236 : v3_1517448501_244;
   assign v3_1517448501_246 = f40 ? v3_1517448501_234 : v3_1517448501_245;
   assign v3_1517448501_247 = f42 ? v3_1517448501_232 : v3_1517448501_246;
   assign v3_1517448501_248 = f44 ? v3_1517448501_230 : v3_1517448501_247;
   assign v3_1517448501_249 = f46 ? v3_1517448501_228 : v3_1517448501_248;
   assign v3_1517448501_250 = f48 ? v3_1517448501_226 : v3_1517448501_249;
   assign v3_1517448501_251 = f50 ? v3_1517448501_224 : v3_1517448501_250;
   assign v3_1517448501_252 = f52 ? v3_1517448501_222 : v3_1517448501_251;
   assign v3_1517448501_253 = f54 ? v3_1517448501_220 : v3_1517448501_252;
   assign v3_1517448501_254 = f56 ? v3_1517448501_218 : v3_1517448501_253;
   assign v3_1517448501_255 = f58 ? v3_1517448501_216 : v3_1517448501_254;
   assign v3_1517448501_256 = f60 ? v3_1517448501_214 : v3_1517448501_255;
   assign v3_1517448501_257 = f62 ? v3_1517448501_212 : v3_1517448501_256;
   assign v3_1517448501_258 = f64 ? v3_1517448501_210 : v3_1517448501_257;
   assign v3_1517448501_259 = f66 ? v3_1517448501_208 : v3_1517448501_258;
   assign v3_1517448501_260 = f68 ? v3_1517448501_206 : v3_1517448501_259;
   assign v3_1517448501_261 = f70 ? v3_1517448501_204 : v3_1517448501_260;
   assign v3_1517448501_262 = f72 ? v3_1517448501_202 : v3_1517448501_261;
   assign v3_1517448501_263 = f74 ? v3_1517448501_200 : v3_1517448501_262;
   assign v3_1517448501_264 = f76 ? v3_1517448501_198 : v3_1517448501_263;
   assign v3_1517448501_265 = f90 ? v3_1517448501_196 : v3_1517448501_264;
   assign v3_1517448501_266 = f93 ? v3_1517448501_187 : v3_1517448501_265;
   assign v3_1517448501_267 = f96 ? v3_1517448501_178 : v3_1517448501_266;
   assign v3_1517448501_268 = 16'b00000000_00000000; 
   assign v3_1517448501_270 = {v_m_responder_0, v3_1517448501_53};
   assign v3_1517448501_271 = v3_1517448501_274 ? ~v3_1517448501_273 : v3_1517448501_272;
   assign v3_1517448501_272 = v3_1517448501_270 >> v3_1517448501_55;
   assign v3_1517448501_273 = ~v3_1517448501_270 >> v3_1517448501_55;
   assign v3_1517448501_274 = v3_1517448501_270[31];
   assign v3_1517448501_275 = v3_1517448501_276 ? v3_1517448501_284 : v3_1517448501_283;
   assign v3_1517448501_276 = v3_1517448501_271[31];
   assign v3_1517448501_277 = v3_1517448501_111[31];
   assign v3_1517448501_278 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_279 = ~v3_1517448501_271 + v3_1517448501_278;
   assign v3_1517448501_280 = ~v3_1517448501_111 + v3_1517448501_278;
   assign v3_1517448501_281 = v3_1517448501_276 ? v3_1517448501_279 : v3_1517448501_271;
   assign v3_1517448501_282 = v3_1517448501_277 ? v3_1517448501_280 : v3_1517448501_111;
   assign v3_1517448501_283 = v3_1517448501_281 % v3_1517448501_282;
   assign v3_1517448501_284 = ~v3_1517448501_283 + v3_1517448501_278;
   assign v3_1517448501_285 = v3_1517448501_288 ? v3_1517448501_295 : v3_1517448501_294;
   assign v3_1517448501_286 = v3_1517448501_275[31];
   assign v3_1517448501_287 = v3_1517448501_77[31];
   assign v3_1517448501_288 = v3_1517448501_286 ^ v3_1517448501_287;
   assign v3_1517448501_289 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_290 = ~v3_1517448501_275 + v3_1517448501_289;
   assign v3_1517448501_291 = ~v3_1517448501_77 + v3_1517448501_289;
   assign v3_1517448501_292 = v3_1517448501_286 ? v3_1517448501_290 : v3_1517448501_275;
   assign v3_1517448501_293 = v3_1517448501_287 ? v3_1517448501_291 : v3_1517448501_77;
   assign v3_1517448501_294 = v3_1517448501_292 / v3_1517448501_293;
   assign v3_1517448501_295 = ~v3_1517448501_294 + v3_1517448501_289;
   assign v3_1517448501_296 = v3_1517448501_285[15:0];
   assign v3_1517448501_297 = f04 ? v3_1517448501_296 : v_party_responder_0;
   assign v3_1517448501_298 = 16'b00000000_00000000; 
   assign v3_1517448501_299 = v3_1517448501_300 ? v3_1517448501_308 : v3_1517448501_307;
   assign v3_1517448501_300 = v3_1517448501_271[31];
   assign v3_1517448501_301 = v3_1517448501_77[31];
   assign v3_1517448501_302 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_303 = ~v3_1517448501_271 + v3_1517448501_302;
   assign v3_1517448501_304 = ~v3_1517448501_77 + v3_1517448501_302;
   assign v3_1517448501_305 = v3_1517448501_300 ? v3_1517448501_303 : v3_1517448501_271;
   assign v3_1517448501_306 = v3_1517448501_301 ? v3_1517448501_304 : v3_1517448501_77;
   assign v3_1517448501_307 = v3_1517448501_305 % v3_1517448501_306;
   assign v3_1517448501_308 = ~v3_1517448501_307 + v3_1517448501_302;
   assign v3_1517448501_309 = v3_1517448501_299[15:0];
   assign v3_1517448501_310 = f04 ? v3_1517448501_309 : v_party_nonce_responder_0;
   assign v3_1517448501_311 = 16'b00000000_00000000; 
   assign v3_1517448501_338 = f31 ? v3_1517448501_208 : v_m_responder_1;
   assign v3_1517448501_339 = f34 ? v3_1517448501_240 : v3_1517448501_338;
   assign v3_1517448501_340 = f37 ? v3_1517448501_238 : v3_1517448501_339;
   assign v3_1517448501_341 = f39 ? v3_1517448501_236 : v3_1517448501_340;
   assign v3_1517448501_342 = f41 ? v3_1517448501_234 : v3_1517448501_341;
   assign v3_1517448501_343 = f43 ? v3_1517448501_232 : v3_1517448501_342;
   assign v3_1517448501_344 = f45 ? v3_1517448501_230 : v3_1517448501_343;
   assign v3_1517448501_345 = f47 ? v3_1517448501_228 : v3_1517448501_344;
   assign v3_1517448501_346 = f49 ? v3_1517448501_226 : v3_1517448501_345;
   assign v3_1517448501_347 = f51 ? v3_1517448501_224 : v3_1517448501_346;
   assign v3_1517448501_348 = f53 ? v3_1517448501_222 : v3_1517448501_347;
   assign v3_1517448501_349 = f55 ? v3_1517448501_220 : v3_1517448501_348;
   assign v3_1517448501_350 = f57 ? v3_1517448501_218 : v3_1517448501_349;
   assign v3_1517448501_351 = f59 ? v3_1517448501_216 : v3_1517448501_350;
   assign v3_1517448501_352 = f61 ? v3_1517448501_214 : v3_1517448501_351;
   assign v3_1517448501_353 = f63 ? v3_1517448501_212 : v3_1517448501_352;
   assign v3_1517448501_354 = f65 ? v3_1517448501_210 : v3_1517448501_353;
   assign v3_1517448501_355 = f67 ? v3_1517448501_208 : v3_1517448501_354;
   assign v3_1517448501_356 = f69 ? v3_1517448501_206 : v3_1517448501_355;
   assign v3_1517448501_357 = f71 ? v3_1517448501_204 : v3_1517448501_356;
   assign v3_1517448501_358 = f73 ? v3_1517448501_202 : v3_1517448501_357;
   assign v3_1517448501_359 = f75 ? v3_1517448501_200 : v3_1517448501_358;
   assign v3_1517448501_360 = f77 ? v3_1517448501_198 : v3_1517448501_359;
   assign v3_1517448501_361 = f91 ? v3_1517448501_196 : v3_1517448501_360;
   assign v3_1517448501_362 = f94 ? v3_1517448501_187 : v3_1517448501_361;
   assign v3_1517448501_363 = f97 ? v3_1517448501_178 : v3_1517448501_362;
   assign v3_1517448501_364 = 16'b00000000_00000000; 
   assign v3_1517448501_366 = {v_m_responder_1, v3_1517448501_53};
   assign v3_1517448501_367 = v3_1517448501_370 ? ~v3_1517448501_369 : v3_1517448501_368;
   assign v3_1517448501_368 = v3_1517448501_366 >> v3_1517448501_55;
   assign v3_1517448501_369 = ~v3_1517448501_366 >> v3_1517448501_55;
   assign v3_1517448501_370 = v3_1517448501_366[31];
   assign v3_1517448501_371 = v3_1517448501_372 ? v3_1517448501_380 : v3_1517448501_379;
   assign v3_1517448501_372 = v3_1517448501_367[31];
   assign v3_1517448501_373 = v3_1517448501_111[31];
   assign v3_1517448501_374 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_375 = ~v3_1517448501_367 + v3_1517448501_374;
   assign v3_1517448501_376 = ~v3_1517448501_111 + v3_1517448501_374;
   assign v3_1517448501_377 = v3_1517448501_372 ? v3_1517448501_375 : v3_1517448501_367;
   assign v3_1517448501_378 = v3_1517448501_373 ? v3_1517448501_376 : v3_1517448501_111;
   assign v3_1517448501_379 = v3_1517448501_377 % v3_1517448501_378;
   assign v3_1517448501_380 = ~v3_1517448501_379 + v3_1517448501_374;
   assign v3_1517448501_381 = v3_1517448501_384 ? v3_1517448501_391 : v3_1517448501_390;
   assign v3_1517448501_382 = v3_1517448501_371[31];
   assign v3_1517448501_383 = v3_1517448501_77[31];
   assign v3_1517448501_384 = v3_1517448501_382 ^ v3_1517448501_383;
   assign v3_1517448501_385 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_386 = ~v3_1517448501_371 + v3_1517448501_385;
   assign v3_1517448501_387 = ~v3_1517448501_77 + v3_1517448501_385;
   assign v3_1517448501_388 = v3_1517448501_382 ? v3_1517448501_386 : v3_1517448501_371;
   assign v3_1517448501_389 = v3_1517448501_383 ? v3_1517448501_387 : v3_1517448501_77;
   assign v3_1517448501_390 = v3_1517448501_388 / v3_1517448501_389;
   assign v3_1517448501_391 = ~v3_1517448501_390 + v3_1517448501_385;
   assign v3_1517448501_392 = v3_1517448501_381[15:0];
   assign v3_1517448501_393 = f08 ? v3_1517448501_392 : v_party_responder_1;
   assign v3_1517448501_394 = 16'b00000000_00000000; 
   assign v3_1517448501_395 = v3_1517448501_396 ? v3_1517448501_404 : v3_1517448501_403;
   assign v3_1517448501_396 = v3_1517448501_367[31];
   assign v3_1517448501_397 = v3_1517448501_77[31];
   assign v3_1517448501_398 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_399 = ~v3_1517448501_367 + v3_1517448501_398;
   assign v3_1517448501_400 = ~v3_1517448501_77 + v3_1517448501_398;
   assign v3_1517448501_401 = v3_1517448501_396 ? v3_1517448501_399 : v3_1517448501_367;
   assign v3_1517448501_402 = v3_1517448501_397 ? v3_1517448501_400 : v3_1517448501_77;
   assign v3_1517448501_403 = v3_1517448501_401 % v3_1517448501_402;
   assign v3_1517448501_404 = ~v3_1517448501_403 + v3_1517448501_398;
   assign v3_1517448501_405 = v3_1517448501_395[15:0];
   assign v3_1517448501_406 = f08 ? v3_1517448501_405 : v_party_nonce_responder_1;
   assign v3_1517448501_407 = 16'b00000000_00000000; 
   assign v3_1517448501_409 = 8'b00000001; 
   assign v3_1517448501_411 = f15 ? v3_1517448501_409 : v_kNa;
   assign v3_1517448501_412 = f25 ? v3_1517448501_409 : v3_1517448501_411;
   assign v3_1517448501_413 = 8'b00000000; 
   assign v3_1517448501_416 = f16 ? v3_1517448501_409 : v_kNb;
   assign v3_1517448501_417 = f26 ? v3_1517448501_409 : v3_1517448501_416;
   assign v3_1517448501_418 = 8'b00000000; 
   assign v3_1517448501_420 = f21 ? v3_1517448501_409 : v_k_Na_Nb__A;
   assign v3_1517448501_421 = 8'b00000000; 
   assign v3_1517448501_423 = f20 ? v3_1517448501_409 : v_k_Na_A__B;
   assign v3_1517448501_424 = 8'b00000000; 
   assign v3_1517448501_427 = f18 ? v3_1517448501_409 : v_k_Nb__B;
   assign v3_1517448501_428 = f28 ? v3_1517448501_409 : v3_1517448501_427;
   assign v3_1517448501_429 = 8'b00000000; 
   assign v3_1517448501_436 = f32 ? v3_1517448501_208 : v_m_intruder;
   assign v3_1517448501_437 = f35 ? v3_1517448501_240 : v3_1517448501_436;
   assign v3_1517448501_438 = f80 ? v3_1517448501_98 : v3_1517448501_437;
   assign v3_1517448501_439 = f83 ? v3_1517448501_86 : v3_1517448501_438;
   assign v3_1517448501_440 = f92 ? v3_1517448501_196 : v3_1517448501_439;
   assign v3_1517448501_441 = f95 ? v3_1517448501_187 : v3_1517448501_440;
   assign v3_1517448501_442 = 16'b00000000_00000000; 
   assign v3_1517448501_443 = ~a_start_initiator_0 & ~f30;
   assign v3_1517448501_444 = v3_1517448501_443 & ~f31;
   assign v3_1517448501_445 = v3_1517448501_444 & ~f32;
   assign v3_1517448501_446 = 1'b0; 
   assign v3_1517448501_447 = ~v3_1517448501_448;
   assign v3_1517448501_448 = ~a_wait_resp_initiator_0 & ~f30;
   assign v3_1517448501_449 = ~v3_1517448501_450;
   assign v3_1517448501_450 = ~v3_1517448501_447 & ~f31;
   assign v3_1517448501_451 = ~v3_1517448501_452;
   assign v3_1517448501_452 = ~v3_1517448501_449 & ~f32;
   assign v3_1517448501_453 = v3_1517448501_451 & ~f78;
   assign v3_1517448501_454 = v3_1517448501_453 & ~f81;
   assign v3_1517448501_455 = v3_1517448501_454 & ~f84;
   assign v3_1517448501_456 = v3_1517448501_455 & ~f86;
   assign v3_1517448501_457 = v3_1517448501_456 & ~f88;
   assign v3_1517448501_458 = 1'b0; 
   assign v3_1517448501_459 = a_got_resp_initiator_0 & ~f00;
   assign v3_1517448501_461 = v3_1517448501_459 & ~f01;
   assign v3_1517448501_462 = ~v3_1517448501_463;
   assign v3_1517448501_463 = ~v3_1517448501_461 & ~f78;
   assign v3_1517448501_464 = ~v3_1517448501_465;
   assign v3_1517448501_465 = ~v3_1517448501_462 & ~f81;
   assign v3_1517448501_466 = ~v3_1517448501_467;
   assign v3_1517448501_467 = ~v3_1517448501_464 & ~f84;
   assign v3_1517448501_468 = ~v3_1517448501_469;
   assign v3_1517448501_469 = ~v3_1517448501_466 & ~f86;
   assign v3_1517448501_470 = ~v3_1517448501_471;
   assign v3_1517448501_471 = ~v3_1517448501_468 & ~f88;
   assign v3_1517448501_472 = 1'b0; 
   assign v3_1517448501_473 = ~v3_1517448501_474;
   assign v3_1517448501_474 = ~a_commited_initiator_0 & ~f00;
   assign v3_1517448501_475 = v3_1517448501_473 & ~f90;
   assign v3_1517448501_476 = v3_1517448501_475 & ~f91;
   assign v3_1517448501_477 = v3_1517448501_476 & ~f92;
   assign v3_1517448501_478 = 1'b0; 
   assign v3_1517448501_479 = ~v3_1517448501_480;
   assign v3_1517448501_480 = ~a_finished_initiator_0 & ~f90;
   assign v3_1517448501_481 = ~v3_1517448501_482;
   assign v3_1517448501_482 = ~v3_1517448501_479 & ~f91;
   assign v3_1517448501_483 = ~v3_1517448501_484;
   assign v3_1517448501_484 = ~v3_1517448501_481 & ~f92;
   assign v3_1517448501_485 = 1'b0; 
   assign v3_1517448501_486 = ~v3_1517448501_487;
   assign v3_1517448501_487 = ~a_corrupted_initiator_0 & ~f01;
   assign v3_1517448501_488 = 1'b0; 
   assign v3_1517448501_489 = ~a_start_initiator_1 & ~f33;
   assign v3_1517448501_490 = v3_1517448501_489 & ~f34;
   assign v3_1517448501_491 = v3_1517448501_490 & ~f35;
   assign v3_1517448501_492 = 1'b0; 
   assign v3_1517448501_493 = ~v3_1517448501_494;
   assign v3_1517448501_494 = ~a_wait_resp_initiator_1 & ~f33;
   assign v3_1517448501_495 = ~v3_1517448501_496;
   assign v3_1517448501_496 = ~v3_1517448501_493 & ~f34;
   assign v3_1517448501_497 = ~v3_1517448501_498;
   assign v3_1517448501_498 = ~v3_1517448501_495 & ~f35;
   assign v3_1517448501_499 = v3_1517448501_497 & ~f79;
   assign v3_1517448501_500 = v3_1517448501_499 & ~f82;
   assign v3_1517448501_501 = v3_1517448501_500 & ~f85;
   assign v3_1517448501_502 = v3_1517448501_501 & ~f87;
   assign v3_1517448501_503 = v3_1517448501_502 & ~f89;
   assign v3_1517448501_504 = 1'b0; 
   assign v3_1517448501_505 = a_got_resp_initiator_1 & ~f02;
   assign v3_1517448501_507 = v3_1517448501_505 & ~f03;
   assign v3_1517448501_508 = ~v3_1517448501_509;
   assign v3_1517448501_509 = ~v3_1517448501_507 & ~f79;
   assign v3_1517448501_510 = ~v3_1517448501_511;
   assign v3_1517448501_511 = ~v3_1517448501_508 & ~f82;
   assign v3_1517448501_512 = ~v3_1517448501_513;
   assign v3_1517448501_513 = ~v3_1517448501_510 & ~f85;
   assign v3_1517448501_514 = ~v3_1517448501_515;
   assign v3_1517448501_515 = ~v3_1517448501_512 & ~f87;
   assign v3_1517448501_516 = ~v3_1517448501_517;
   assign v3_1517448501_517 = ~v3_1517448501_514 & ~f89;
   assign v3_1517448501_518 = 1'b0; 
   assign v3_1517448501_519 = ~v3_1517448501_520;
   assign v3_1517448501_520 = ~a_commited_initiator_1 & ~f02;
   assign v3_1517448501_521 = v3_1517448501_519 & ~f93;
   assign v3_1517448501_522 = v3_1517448501_521 & ~f94;
   assign v3_1517448501_523 = v3_1517448501_522 & ~f95;
   assign v3_1517448501_524 = 1'b0; 
   assign v3_1517448501_525 = ~v3_1517448501_526;
   assign v3_1517448501_526 = ~a_finished_initiator_1 & ~f93;
   assign v3_1517448501_527 = ~v3_1517448501_528;
   assign v3_1517448501_528 = ~v3_1517448501_525 & ~f94;
   assign v3_1517448501_529 = ~v3_1517448501_530;
   assign v3_1517448501_530 = ~v3_1517448501_527 & ~f95;
   assign v3_1517448501_531 = 1'b0; 
   assign v3_1517448501_532 = ~v3_1517448501_533;
   assign v3_1517448501_533 = ~a_corrupted_initiator_1 & ~f03;
   assign v3_1517448501_534 = 1'b0; 
   assign v3_1517448501_535 = ~a_start_responder_0 & ~f30;
   assign v3_1517448501_536 = v3_1517448501_535 & ~f33;
   assign v3_1517448501_537 = v3_1517448501_536 & ~f36;
   assign v3_1517448501_538 = v3_1517448501_537 & ~f38;
   assign v3_1517448501_539 = v3_1517448501_538 & ~f40;
   assign v3_1517448501_540 = v3_1517448501_539 & ~f42;
   assign v3_1517448501_541 = v3_1517448501_540 & ~f44;
   assign v3_1517448501_542 = v3_1517448501_541 & ~f46;
   assign v3_1517448501_543 = v3_1517448501_542 & ~f48;
   assign v3_1517448501_544 = v3_1517448501_543 & ~f50;
   assign v3_1517448501_545 = v3_1517448501_544 & ~f52;
   assign v3_1517448501_546 = v3_1517448501_545 & ~f54;
   assign v3_1517448501_547 = v3_1517448501_546 & ~f56;
   assign v3_1517448501_548 = v3_1517448501_547 & ~f58;
   assign v3_1517448501_549 = v3_1517448501_548 & ~f60;
   assign v3_1517448501_550 = v3_1517448501_549 & ~f62;
   assign v3_1517448501_551 = v3_1517448501_550 & ~f64;
   assign v3_1517448501_552 = v3_1517448501_551 & ~f66;
   assign v3_1517448501_553 = v3_1517448501_552 & ~f68;
   assign v3_1517448501_554 = v3_1517448501_553 & ~f70;
   assign v3_1517448501_555 = v3_1517448501_554 & ~f72;
   assign v3_1517448501_556 = v3_1517448501_555 & ~f74;
   assign v3_1517448501_557 = v3_1517448501_556 & ~f76;
   assign v3_1517448501_558 = 1'b0; 
   assign v3_1517448501_559 = a_got_msg_responder_0 & ~f04;
   assign v3_1517448501_561 = v3_1517448501_559 & ~f05;
   assign v3_1517448501_562 = ~v3_1517448501_563;
   assign v3_1517448501_563 = ~v3_1517448501_561 & ~f30;
   assign v3_1517448501_564 = ~v3_1517448501_565;
   assign v3_1517448501_565 = ~v3_1517448501_562 & ~f33;
   assign v3_1517448501_566 = ~v3_1517448501_567;
   assign v3_1517448501_567 = ~v3_1517448501_564 & ~f36;
   assign v3_1517448501_568 = ~v3_1517448501_569;
   assign v3_1517448501_569 = ~v3_1517448501_566 & ~f38;
   assign v3_1517448501_570 = ~v3_1517448501_571;
   assign v3_1517448501_571 = ~v3_1517448501_568 & ~f40;
   assign v3_1517448501_572 = ~v3_1517448501_573;
   assign v3_1517448501_573 = ~v3_1517448501_570 & ~f42;
   assign v3_1517448501_574 = ~v3_1517448501_575;
   assign v3_1517448501_575 = ~v3_1517448501_572 & ~f44;
   assign v3_1517448501_576 = ~v3_1517448501_577;
   assign v3_1517448501_577 = ~v3_1517448501_574 & ~f46;
   assign v3_1517448501_578 = ~v3_1517448501_579;
   assign v3_1517448501_579 = ~v3_1517448501_576 & ~f48;
   assign v3_1517448501_580 = ~v3_1517448501_581;
   assign v3_1517448501_581 = ~v3_1517448501_578 & ~f50;
   assign v3_1517448501_582 = ~v3_1517448501_583;
   assign v3_1517448501_583 = ~v3_1517448501_580 & ~f52;
   assign v3_1517448501_584 = ~v3_1517448501_585;
   assign v3_1517448501_585 = ~v3_1517448501_582 & ~f54;
   assign v3_1517448501_586 = ~v3_1517448501_587;
   assign v3_1517448501_587 = ~v3_1517448501_584 & ~f56;
   assign v3_1517448501_588 = ~v3_1517448501_589;
   assign v3_1517448501_589 = ~v3_1517448501_586 & ~f58;
   assign v3_1517448501_590 = ~v3_1517448501_591;
   assign v3_1517448501_591 = ~v3_1517448501_588 & ~f60;
   assign v3_1517448501_592 = ~v3_1517448501_593;
   assign v3_1517448501_593 = ~v3_1517448501_590 & ~f62;
   assign v3_1517448501_594 = ~v3_1517448501_595;
   assign v3_1517448501_595 = ~v3_1517448501_592 & ~f64;
   assign v3_1517448501_596 = ~v3_1517448501_597;
   assign v3_1517448501_597 = ~v3_1517448501_594 & ~f66;
   assign v3_1517448501_598 = ~v3_1517448501_599;
   assign v3_1517448501_599 = ~v3_1517448501_596 & ~f68;
   assign v3_1517448501_600 = ~v3_1517448501_601;
   assign v3_1517448501_601 = ~v3_1517448501_598 & ~f70;
   assign v3_1517448501_602 = ~v3_1517448501_603;
   assign v3_1517448501_603 = ~v3_1517448501_600 & ~f72;
   assign v3_1517448501_604 = ~v3_1517448501_605;
   assign v3_1517448501_605 = ~v3_1517448501_602 & ~f74;
   assign v3_1517448501_606 = ~v3_1517448501_607;
   assign v3_1517448501_607 = ~v3_1517448501_604 & ~f76;
   assign v3_1517448501_608 = 1'b0; 
   assign v3_1517448501_609 = ~v3_1517448501_610;
   assign v3_1517448501_610 = ~a_send_reply_responder_0 & ~f04;
   assign v3_1517448501_611 = v3_1517448501_609 & ~f78;
   assign v3_1517448501_612 = v3_1517448501_611 & ~f79;
   assign v3_1517448501_613 = v3_1517448501_612 & ~f80;
   assign v3_1517448501_614 = 1'b0; 
   assign v3_1517448501_615 = ~v3_1517448501_616;
   assign v3_1517448501_616 = ~a_wait_resp_responder_0 & ~f78;
   assign v3_1517448501_617 = ~v3_1517448501_618;
   assign v3_1517448501_618 = ~v3_1517448501_615 & ~f79;
   assign v3_1517448501_619 = ~v3_1517448501_620;
   assign v3_1517448501_620 = ~v3_1517448501_617 & ~f80;
   assign v3_1517448501_621 = v3_1517448501_619 & ~f90;
   assign v3_1517448501_622 = v3_1517448501_621 & ~f93;
   assign v3_1517448501_623 = v3_1517448501_622 & ~f96;
   assign v3_1517448501_624 = 1'b0; 
   assign v3_1517448501_626 = a_got_resp_responder_0 & ~f06;
   assign v3_1517448501_628 = v3_1517448501_626 & ~f07;
   assign v3_1517448501_629 = ~v3_1517448501_630;
   assign v3_1517448501_630 = ~v3_1517448501_628 & ~f90;
   assign v3_1517448501_631 = ~v3_1517448501_632;
   assign v3_1517448501_632 = ~v3_1517448501_629 & ~f93;
   assign v3_1517448501_633 = ~v3_1517448501_634;
   assign v3_1517448501_634 = ~v3_1517448501_631 & ~f96;
   assign v3_1517448501_635 = 1'b0; 
   assign v3_1517448501_636 = ~v3_1517448501_637;
   assign v3_1517448501_637 = ~a_finished_responder_0 & ~f07;
   assign v3_1517448501_638 = 1'b0; 
   assign v3_1517448501_639 = ~v3_1517448501_640;
   assign v3_1517448501_640 = ~a_corrupted_responder_0 & ~f05;
   assign v3_1517448501_641 = ~v3_1517448501_642;
   assign v3_1517448501_642 = ~v3_1517448501_639 & ~f06;
   assign v3_1517448501_643 = 1'b0; 
   assign v3_1517448501_644 = ~a_start_responder_1 & ~f31;
   assign v3_1517448501_645 = v3_1517448501_644 & ~f34;
   assign v3_1517448501_646 = v3_1517448501_645 & ~f37;
   assign v3_1517448501_647 = v3_1517448501_646 & ~f39;
   assign v3_1517448501_648 = v3_1517448501_647 & ~f41;
   assign v3_1517448501_649 = v3_1517448501_648 & ~f43;
   assign v3_1517448501_650 = v3_1517448501_649 & ~f45;
   assign v3_1517448501_651 = v3_1517448501_650 & ~f47;
   assign v3_1517448501_652 = v3_1517448501_651 & ~f49;
   assign v3_1517448501_653 = v3_1517448501_652 & ~f51;
   assign v3_1517448501_654 = v3_1517448501_653 & ~f53;
   assign v3_1517448501_655 = v3_1517448501_654 & ~f55;
   assign v3_1517448501_656 = v3_1517448501_655 & ~f57;
   assign v3_1517448501_657 = v3_1517448501_656 & ~f59;
   assign v3_1517448501_658 = v3_1517448501_657 & ~f61;
   assign v3_1517448501_659 = v3_1517448501_658 & ~f63;
   assign v3_1517448501_660 = v3_1517448501_659 & ~f65;
   assign v3_1517448501_661 = v3_1517448501_660 & ~f67;
   assign v3_1517448501_662 = v3_1517448501_661 & ~f69;
   assign v3_1517448501_663 = v3_1517448501_662 & ~f71;
   assign v3_1517448501_664 = v3_1517448501_663 & ~f73;
   assign v3_1517448501_665 = v3_1517448501_664 & ~f75;
   assign v3_1517448501_666 = v3_1517448501_665 & ~f77;
   assign v3_1517448501_667 = 1'b0; 
   assign v3_1517448501_668 = a_got_msg_responder_1 & ~f08;
   assign v3_1517448501_670 = v3_1517448501_668 & ~f09;
   assign v3_1517448501_671 = ~v3_1517448501_672;
   assign v3_1517448501_672 = ~v3_1517448501_670 & ~f31;
   assign v3_1517448501_673 = ~v3_1517448501_674;
   assign v3_1517448501_674 = ~v3_1517448501_671 & ~f34;
   assign v3_1517448501_675 = ~v3_1517448501_676;
   assign v3_1517448501_676 = ~v3_1517448501_673 & ~f37;
   assign v3_1517448501_677 = ~v3_1517448501_678;
   assign v3_1517448501_678 = ~v3_1517448501_675 & ~f39;
   assign v3_1517448501_679 = ~v3_1517448501_680;
   assign v3_1517448501_680 = ~v3_1517448501_677 & ~f41;
   assign v3_1517448501_681 = ~v3_1517448501_682;
   assign v3_1517448501_682 = ~v3_1517448501_679 & ~f43;
   assign v3_1517448501_683 = ~v3_1517448501_684;
   assign v3_1517448501_684 = ~v3_1517448501_681 & ~f45;
   assign v3_1517448501_685 = ~v3_1517448501_686;
   assign v3_1517448501_686 = ~v3_1517448501_683 & ~f47;
   assign v3_1517448501_687 = ~v3_1517448501_688;
   assign v3_1517448501_688 = ~v3_1517448501_685 & ~f49;
   assign v3_1517448501_689 = ~v3_1517448501_690;
   assign v3_1517448501_690 = ~v3_1517448501_687 & ~f51;
   assign v3_1517448501_691 = ~v3_1517448501_692;
   assign v3_1517448501_692 = ~v3_1517448501_689 & ~f53;
   assign v3_1517448501_693 = ~v3_1517448501_694;
   assign v3_1517448501_694 = ~v3_1517448501_691 & ~f55;
   assign v3_1517448501_695 = ~v3_1517448501_696;
   assign v3_1517448501_696 = ~v3_1517448501_693 & ~f57;
   assign v3_1517448501_697 = ~v3_1517448501_698;
   assign v3_1517448501_698 = ~v3_1517448501_695 & ~f59;
   assign v3_1517448501_699 = ~v3_1517448501_700;
   assign v3_1517448501_700 = ~v3_1517448501_697 & ~f61;
   assign v3_1517448501_701 = ~v3_1517448501_702;
   assign v3_1517448501_702 = ~v3_1517448501_699 & ~f63;
   assign v3_1517448501_703 = ~v3_1517448501_704;
   assign v3_1517448501_704 = ~v3_1517448501_701 & ~f65;
   assign v3_1517448501_705 = ~v3_1517448501_706;
   assign v3_1517448501_706 = ~v3_1517448501_703 & ~f67;
   assign v3_1517448501_707 = ~v3_1517448501_708;
   assign v3_1517448501_708 = ~v3_1517448501_705 & ~f69;
   assign v3_1517448501_709 = ~v3_1517448501_710;
   assign v3_1517448501_710 = ~v3_1517448501_707 & ~f71;
   assign v3_1517448501_711 = ~v3_1517448501_712;
   assign v3_1517448501_712 = ~v3_1517448501_709 & ~f73;
   assign v3_1517448501_713 = ~v3_1517448501_714;
   assign v3_1517448501_714 = ~v3_1517448501_711 & ~f75;
   assign v3_1517448501_715 = ~v3_1517448501_716;
   assign v3_1517448501_716 = ~v3_1517448501_713 & ~f77;
   assign v3_1517448501_717 = 1'b0; 
   assign v3_1517448501_718 = ~v3_1517448501_719;
   assign v3_1517448501_719 = ~a_send_reply_responder_1 & ~f08;
   assign v3_1517448501_720 = v3_1517448501_718 & ~f81;
   assign v3_1517448501_721 = v3_1517448501_720 & ~f82;
   assign v3_1517448501_722 = v3_1517448501_721 & ~f83;
   assign v3_1517448501_723 = 1'b0; 
   assign v3_1517448501_724 = ~v3_1517448501_725;
   assign v3_1517448501_725 = ~a_wait_resp_responder_1 & ~f81;
   assign v3_1517448501_726 = ~v3_1517448501_727;
   assign v3_1517448501_727 = ~v3_1517448501_724 & ~f82;
   assign v3_1517448501_728 = ~v3_1517448501_729;
   assign v3_1517448501_729 = ~v3_1517448501_726 & ~f83;
   assign v3_1517448501_730 = v3_1517448501_728 & ~f91;
   assign v3_1517448501_731 = v3_1517448501_730 & ~f94;
   assign v3_1517448501_732 = v3_1517448501_731 & ~f97;
   assign v3_1517448501_733 = 1'b0; 
   assign v3_1517448501_735 = a_got_resp_responder_1 & ~f10;
   assign v3_1517448501_737 = v3_1517448501_735 & ~f11;
   assign v3_1517448501_738 = ~v3_1517448501_739;
   assign v3_1517448501_739 = ~v3_1517448501_737 & ~f91;
   assign v3_1517448501_740 = ~v3_1517448501_741;
   assign v3_1517448501_741 = ~v3_1517448501_738 & ~f94;
   assign v3_1517448501_742 = ~v3_1517448501_743;
   assign v3_1517448501_743 = ~v3_1517448501_740 & ~f97;
   assign v3_1517448501_744 = 1'b0; 
   assign v3_1517448501_745 = ~v3_1517448501_746;
   assign v3_1517448501_746 = ~a_finished_responder_1 & ~f11;
   assign v3_1517448501_747 = 1'b0; 
   assign v3_1517448501_748 = ~v3_1517448501_749;
   assign v3_1517448501_749 = ~a_corrupted_responder_1 & ~f09;
   assign v3_1517448501_750 = ~v3_1517448501_751;
   assign v3_1517448501_751 = ~v3_1517448501_748 & ~f10;
   assign v3_1517448501_752 = 1'b0; 
   assign v3_1517448501_754 = ~v3_1517448501_755;
   assign v3_1517448501_755 = a_q & ~f12;
   assign v3_1517448501_756 = ~v3_1517448501_757;
   assign v3_1517448501_757 = ~v3_1517448501_754 & ~f18;
   assign v3_1517448501_759 = ~v3_1517448501_760;
   assign v3_1517448501_760 = ~v3_1517448501_756 & ~f19;
   assign v3_1517448501_761 = ~v3_1517448501_762;
   assign v3_1517448501_762 = ~v3_1517448501_759 & ~f20;
   assign v3_1517448501_763 = ~v3_1517448501_764;
   assign v3_1517448501_764 = ~v3_1517448501_761 & ~f21;
   assign v3_1517448501_766 = ~v3_1517448501_767;
   assign v3_1517448501_767 = ~v3_1517448501_763 & ~f22;
   assign v3_1517448501_768 = ~v3_1517448501_769;
   assign v3_1517448501_769 = ~v3_1517448501_766 & ~f25;
   assign v3_1517448501_770 = ~v3_1517448501_771;
   assign v3_1517448501_771 = ~v3_1517448501_768 & ~f26;
   assign v3_1517448501_773 = ~v3_1517448501_774;
   assign v3_1517448501_774 = ~v3_1517448501_770 & ~f27;
   assign v3_1517448501_775 = ~v3_1517448501_776;
   assign v3_1517448501_776 = ~v3_1517448501_773 & ~f28;
   assign v3_1517448501_778 = ~v3_1517448501_779;
   assign v3_1517448501_779 = ~v3_1517448501_775 & ~f29;
   assign v3_1517448501_780 = v3_1517448501_778 & ~f32;
   assign v3_1517448501_781 = v3_1517448501_780 & ~f35;
   assign v3_1517448501_782 = v3_1517448501_781 & ~f80;
   assign v3_1517448501_783 = v3_1517448501_782 & ~f83;
   assign v3_1517448501_784 = v3_1517448501_783 & ~f92;
   assign v3_1517448501_785 = v3_1517448501_784 & ~f95;
   assign v3_1517448501_786 = 1'b0; 
   assign v3_1517448501_787 = a_got3 & ~f12;
   assign v3_1517448501_789 = v3_1517448501_787 & ~f13;
   assign v3_1517448501_791 = v3_1517448501_789 & ~f14;
   assign v3_1517448501_792 = ~v3_1517448501_793;
   assign v3_1517448501_793 = ~v3_1517448501_791 & ~f32;
   assign v3_1517448501_794 = ~v3_1517448501_795;
   assign v3_1517448501_795 = ~v3_1517448501_792 & ~f35;
   assign v3_1517448501_796 = ~v3_1517448501_797;
   assign v3_1517448501_797 = ~v3_1517448501_794 & ~f80;
   assign v3_1517448501_798 = ~v3_1517448501_799;
   assign v3_1517448501_799 = ~v3_1517448501_796 & ~f83;
   assign v3_1517448501_800 = 1'b0; 
   assign v3_1517448501_801 = ~v3_1517448501_802;
   assign v3_1517448501_802 = ~a_c1 & ~f13;
   assign v3_1517448501_803 = v3_1517448501_801 & ~f15;
   assign v3_1517448501_804 = v3_1517448501_803 & ~f16;
   assign v3_1517448501_806 = v3_1517448501_804 & ~f17;
   assign v3_1517448501_807 = 1'b0; 
   assign v3_1517448501_808 = ~v3_1517448501_809;
   assign v3_1517448501_809 = ~a_c2 & ~f15;
   assign v3_1517448501_810 = ~v3_1517448501_811;
   assign v3_1517448501_811 = ~v3_1517448501_808 & ~f16;
   assign v3_1517448501_812 = ~v3_1517448501_813;
   assign v3_1517448501_813 = ~v3_1517448501_810 & ~f17;
   assign v3_1517448501_814 = v3_1517448501_812 & ~f18;
   assign v3_1517448501_815 = v3_1517448501_814 & ~f19;
   assign v3_1517448501_816 = 1'b0; 
   assign v3_1517448501_817 = ~v3_1517448501_818;
   assign v3_1517448501_818 = ~a_d1 & ~f14;
   assign v3_1517448501_819 = v3_1517448501_817 & ~f20;
   assign v3_1517448501_820 = v3_1517448501_819 & ~f21;
   assign v3_1517448501_821 = v3_1517448501_820 & ~f22;
   assign v3_1517448501_822 = 1'b0; 
   assign v3_1517448501_824 = a_got2 & ~f23;
   assign v3_1517448501_826 = v3_1517448501_824 & ~f24;
   assign v3_1517448501_827 = ~v3_1517448501_828;
   assign v3_1517448501_828 = ~v3_1517448501_826 & ~f92;
   assign v3_1517448501_829 = ~v3_1517448501_830;
   assign v3_1517448501_830 = ~v3_1517448501_827 & ~f95;
   assign v3_1517448501_831 = 1'b0; 
   assign v3_1517448501_832 = ~v3_1517448501_833;
   assign v3_1517448501_833 = ~a_e1 & ~f23;
   assign v3_1517448501_834 = v3_1517448501_832 & ~f25;
   assign v3_1517448501_835 = v3_1517448501_834 & ~f26;
   assign v3_1517448501_836 = v3_1517448501_835 & ~f27;
   assign v3_1517448501_837 = 1'b0; 
   assign v3_1517448501_838 = ~v3_1517448501_839;
   assign v3_1517448501_839 = ~a_f1 & ~f24;
   assign v3_1517448501_840 = v3_1517448501_838 & ~f28;
   assign v3_1517448501_841 = v3_1517448501_840 & ~f29;
   assign v3_1517448501_842 = 1'b0; 
   assign v3_1517448501_843 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_844 = v3_1517448501_845 ? v3_1517448501_853 : v3_1517448501_852;
   assign v3_1517448501_845 = v3_1517448501_107[31];
   assign v3_1517448501_846 = v3_1517448501_77[31];
   assign v3_1517448501_847 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_848 = ~v3_1517448501_107 + v3_1517448501_847;
   assign v3_1517448501_849 = ~v3_1517448501_77 + v3_1517448501_847;
   assign v3_1517448501_850 = v3_1517448501_845 ? v3_1517448501_848 : v3_1517448501_107;
   assign v3_1517448501_851 = v3_1517448501_846 ? v3_1517448501_849 : v3_1517448501_77;
   assign v3_1517448501_852 = v3_1517448501_850 % v3_1517448501_851;
   assign v3_1517448501_853 = ~v3_1517448501_852 + v3_1517448501_847;
   assign v3_1517448501_854 = v3_1517448501_843 == v3_1517448501_844;
   assign v3_1517448501_855 = v3_1517448501_858 ? v3_1517448501_865 : v3_1517448501_864;
   assign v3_1517448501_856 = v3_1517448501_107[31];
   assign v3_1517448501_857 = v3_1517448501_111[31];
   assign v3_1517448501_858 = v3_1517448501_856 ^ v3_1517448501_857;
   assign v3_1517448501_859 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_860 = ~v3_1517448501_107 + v3_1517448501_859;
   assign v3_1517448501_861 = ~v3_1517448501_111 + v3_1517448501_859;
   assign v3_1517448501_862 = v3_1517448501_856 ? v3_1517448501_860 : v3_1517448501_107;
   assign v3_1517448501_863 = v3_1517448501_857 ? v3_1517448501_861 : v3_1517448501_111;
   assign v3_1517448501_864 = v3_1517448501_862 / v3_1517448501_863;
   assign v3_1517448501_865 = ~v3_1517448501_864 + v3_1517448501_859;
   assign v3_1517448501_866 = v3_1517448501_52 == v3_1517448501_855;
   assign v3_1517448501_867 = v3_1517448501_854 & v3_1517448501_866;
   assign v3_1517448501_868 = a_got_resp_initiator_0 & v3_1517448501_867;
   assign v3_1517448501_869 = ~v3_1517448501_870;
   assign v3_1517448501_870 = f00 & ~v3_1517448501_868;
   assign v3_1517448501_871 = a_got_resp_initiator_0 & ~v3_1517448501_867;
   assign v3_1517448501_872 = ~v3_1517448501_873;
   assign v3_1517448501_873 = f01 & ~v3_1517448501_871;
   assign v3_1517448501_874 = v3_1517448501_869 & v3_1517448501_872;
   assign v3_1517448501_875 = 32'b00000000_00000000_00000000_00000010; 
   assign v3_1517448501_876 = v3_1517448501_877 ? v3_1517448501_885 : v3_1517448501_884;
   assign v3_1517448501_877 = v3_1517448501_149[31];
   assign v3_1517448501_878 = v3_1517448501_77[31];
   assign v3_1517448501_879 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_880 = ~v3_1517448501_149 + v3_1517448501_879;
   assign v3_1517448501_881 = ~v3_1517448501_77 + v3_1517448501_879;
   assign v3_1517448501_882 = v3_1517448501_877 ? v3_1517448501_880 : v3_1517448501_149;
   assign v3_1517448501_883 = v3_1517448501_878 ? v3_1517448501_881 : v3_1517448501_77;
   assign v3_1517448501_884 = v3_1517448501_882 % v3_1517448501_883;
   assign v3_1517448501_885 = ~v3_1517448501_884 + v3_1517448501_879;
   assign v3_1517448501_886 = v3_1517448501_875 == v3_1517448501_876;
   assign v3_1517448501_887 = 32'b00000000_00000000_00000000_00001000; 
   assign v3_1517448501_888 = v3_1517448501_891 ? v3_1517448501_898 : v3_1517448501_897;
   assign v3_1517448501_889 = v3_1517448501_149[31];
   assign v3_1517448501_890 = v3_1517448501_111[31];
   assign v3_1517448501_891 = v3_1517448501_889 ^ v3_1517448501_890;
   assign v3_1517448501_892 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_893 = ~v3_1517448501_149 + v3_1517448501_892;
   assign v3_1517448501_894 = ~v3_1517448501_111 + v3_1517448501_892;
   assign v3_1517448501_895 = v3_1517448501_889 ? v3_1517448501_893 : v3_1517448501_149;
   assign v3_1517448501_896 = v3_1517448501_890 ? v3_1517448501_894 : v3_1517448501_111;
   assign v3_1517448501_897 = v3_1517448501_895 / v3_1517448501_896;
   assign v3_1517448501_898 = ~v3_1517448501_897 + v3_1517448501_892;
   assign v3_1517448501_899 = v3_1517448501_887 == v3_1517448501_888;
   assign v3_1517448501_900 = v3_1517448501_886 & v3_1517448501_899;
   assign v3_1517448501_901 = a_got_resp_initiator_1 & v3_1517448501_900;
   assign v3_1517448501_902 = ~v3_1517448501_903;
   assign v3_1517448501_903 = f02 & ~v3_1517448501_901;
   assign v3_1517448501_904 = v3_1517448501_874 & v3_1517448501_902;
   assign v3_1517448501_905 = a_got_resp_initiator_1 & ~v3_1517448501_900;
   assign v3_1517448501_906 = ~v3_1517448501_907;
   assign v3_1517448501_907 = f03 & ~v3_1517448501_905;
   assign v3_1517448501_908 = v3_1517448501_904 & v3_1517448501_906;
   assign v3_1517448501_909 = 32'b00000000_00000000_00000000_00001010; 
   assign v3_1517448501_910 = v3_1517448501_913 ? v3_1517448501_920 : v3_1517448501_919;
   assign v3_1517448501_911 = v3_1517448501_271[31];
   assign v3_1517448501_912 = v3_1517448501_111[31];
   assign v3_1517448501_913 = v3_1517448501_911 ^ v3_1517448501_912;
   assign v3_1517448501_914 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_915 = ~v3_1517448501_271 + v3_1517448501_914;
   assign v3_1517448501_916 = ~v3_1517448501_111 + v3_1517448501_914;
   assign v3_1517448501_917 = v3_1517448501_911 ? v3_1517448501_915 : v3_1517448501_271;
   assign v3_1517448501_918 = v3_1517448501_912 ? v3_1517448501_916 : v3_1517448501_111;
   assign v3_1517448501_919 = v3_1517448501_917 / v3_1517448501_918;
   assign v3_1517448501_920 = ~v3_1517448501_919 + v3_1517448501_914;
   assign v3_1517448501_921 = v3_1517448501_909 == v3_1517448501_910;
   assign v3_1517448501_922 = a_got_msg_responder_0 & v3_1517448501_921;
   assign v3_1517448501_923 = ~v3_1517448501_924;
   assign v3_1517448501_924 = f04 & ~v3_1517448501_922;
   assign v3_1517448501_925 = v3_1517448501_908 & v3_1517448501_923;
   assign v3_1517448501_926 = a_got_msg_responder_0 & ~v3_1517448501_921;
   assign v3_1517448501_927 = ~v3_1517448501_928;
   assign v3_1517448501_928 = f05 & ~v3_1517448501_926;
   assign v3_1517448501_929 = v3_1517448501_925 & v3_1517448501_927;
   assign v3_1517448501_930 = 32'b00000000_00000000_00000000_00000100; 
   assign v3_1517448501_931 = v3_1517448501_930 == v3_1517448501_299;
   assign v3_1517448501_932 = v3_1517448501_909 == v3_1517448501_285;
   assign v3_1517448501_933 = v3_1517448501_931 & v3_1517448501_932;
   assign v3_1517448501_934 = a_got_resp_responder_0 & ~v3_1517448501_933;
   assign v3_1517448501_935 = ~v3_1517448501_936;
   assign v3_1517448501_936 = f06 & ~v3_1517448501_934;
   assign v3_1517448501_937 = v3_1517448501_929 & v3_1517448501_935;
   assign v3_1517448501_938 = a_got_resp_responder_0 & v3_1517448501_933;
   assign v3_1517448501_939 = ~v3_1517448501_940;
   assign v3_1517448501_940 = f07 & ~v3_1517448501_938;
   assign v3_1517448501_941 = v3_1517448501_937 & v3_1517448501_939;
   assign v3_1517448501_942 = 32'b00000000_00000000_00000000_00001011; 
   assign v3_1517448501_943 = v3_1517448501_946 ? v3_1517448501_953 : v3_1517448501_952;
   assign v3_1517448501_944 = v3_1517448501_367[31];
   assign v3_1517448501_945 = v3_1517448501_111[31];
   assign v3_1517448501_946 = v3_1517448501_944 ^ v3_1517448501_945;
   assign v3_1517448501_947 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_948 = ~v3_1517448501_367 + v3_1517448501_947;
   assign v3_1517448501_949 = ~v3_1517448501_111 + v3_1517448501_947;
   assign v3_1517448501_950 = v3_1517448501_944 ? v3_1517448501_948 : v3_1517448501_367;
   assign v3_1517448501_951 = v3_1517448501_945 ? v3_1517448501_949 : v3_1517448501_111;
   assign v3_1517448501_952 = v3_1517448501_950 / v3_1517448501_951;
   assign v3_1517448501_953 = ~v3_1517448501_952 + v3_1517448501_947;
   assign v3_1517448501_954 = v3_1517448501_942 == v3_1517448501_943;
   assign v3_1517448501_955 = a_got_msg_responder_1 & v3_1517448501_954;
   assign v3_1517448501_956 = ~v3_1517448501_957;
   assign v3_1517448501_957 = f08 & ~v3_1517448501_955;
   assign v3_1517448501_958 = v3_1517448501_941 & v3_1517448501_956;
   assign v3_1517448501_959 = a_got_msg_responder_1 & ~v3_1517448501_954;
   assign v3_1517448501_960 = ~v3_1517448501_961;
   assign v3_1517448501_961 = f09 & ~v3_1517448501_959;
   assign v3_1517448501_962 = v3_1517448501_958 & v3_1517448501_960;
   assign v3_1517448501_963 = 32'b00000000_00000000_00000000_00000101; 
   assign v3_1517448501_964 = v3_1517448501_963 == v3_1517448501_395;
   assign v3_1517448501_965 = v3_1517448501_942 == v3_1517448501_381;
   assign v3_1517448501_966 = v3_1517448501_964 & v3_1517448501_965;
   assign v3_1517448501_967 = a_got_resp_responder_1 & ~v3_1517448501_966;
   assign v3_1517448501_968 = ~v3_1517448501_969;
   assign v3_1517448501_969 = f10 & ~v3_1517448501_967;
   assign v3_1517448501_970 = v3_1517448501_962 & v3_1517448501_968;
   assign v3_1517448501_971 = a_got_resp_responder_1 & v3_1517448501_966;
   assign v3_1517448501_972 = ~v3_1517448501_973;
   assign v3_1517448501_973 = f11 & ~v3_1517448501_971;
   assign v3_1517448501_974 = v3_1517448501_970 & v3_1517448501_972;
   assign v3_1517448501_975 = ~v3_1517448501_976;
   assign v3_1517448501_976 = ~a_got3 & f12;
   assign v3_1517448501_977 = v3_1517448501_974 & v3_1517448501_975;
   assign v3_1517448501_978 = {v_m_intruder, v3_1517448501_53};
   assign v3_1517448501_979 = v3_1517448501_982 ? ~v3_1517448501_981 : v3_1517448501_980;
   assign v3_1517448501_980 = v3_1517448501_978 >> v3_1517448501_55;
   assign v3_1517448501_981 = ~v3_1517448501_978 >> v3_1517448501_55;
   assign v3_1517448501_982 = v3_1517448501_978[31];
   assign v3_1517448501_983 = v3_1517448501_986 ? v3_1517448501_993 : v3_1517448501_992;
   assign v3_1517448501_984 = v3_1517448501_979[31];
   assign v3_1517448501_985 = v3_1517448501_111[31];
   assign v3_1517448501_986 = v3_1517448501_984 ^ v3_1517448501_985;
   assign v3_1517448501_987 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_988 = ~v3_1517448501_979 + v3_1517448501_987;
   assign v3_1517448501_989 = ~v3_1517448501_111 + v3_1517448501_987;
   assign v3_1517448501_990 = v3_1517448501_984 ? v3_1517448501_988 : v3_1517448501_979;
   assign v3_1517448501_991 = v3_1517448501_985 ? v3_1517448501_989 : v3_1517448501_111;
   assign v3_1517448501_992 = v3_1517448501_990 / v3_1517448501_991;
   assign v3_1517448501_993 = ~v3_1517448501_992 + v3_1517448501_987;
   assign v3_1517448501_994 = v3_1517448501_875 == v3_1517448501_983;
   assign v3_1517448501_995 = a_got3 & v3_1517448501_994;
   assign v3_1517448501_996 = ~v3_1517448501_997;
   assign v3_1517448501_997 = f13 & ~v3_1517448501_995;
   assign v3_1517448501_998 = v3_1517448501_977 & v3_1517448501_996;
   assign v3_1517448501_999 = a_got3 & ~v3_1517448501_994;
   assign v3_1517448501_1000 = ~v3_1517448501_1001;
   assign v3_1517448501_1001 = f14 & ~v3_1517448501_999;
   assign v3_1517448501_1002 = v3_1517448501_998 & v3_1517448501_1000;
   assign v3_1517448501_1003 = v3_1517448501_1004 ? v3_1517448501_1012 : v3_1517448501_1011;
   assign v3_1517448501_1004 = v3_1517448501_979[31];
   assign v3_1517448501_1005 = v3_1517448501_77[31];
   assign v3_1517448501_1006 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1007 = ~v3_1517448501_979 + v3_1517448501_1006;
   assign v3_1517448501_1008 = ~v3_1517448501_77 + v3_1517448501_1006;
   assign v3_1517448501_1009 = v3_1517448501_1004 ? v3_1517448501_1007 : v3_1517448501_979;
   assign v3_1517448501_1010 = v3_1517448501_1005 ? v3_1517448501_1008 : v3_1517448501_77;
   assign v3_1517448501_1011 = v3_1517448501_1009 % v3_1517448501_1010;
   assign v3_1517448501_1012 = ~v3_1517448501_1011 + v3_1517448501_1006;
   assign v3_1517448501_1013 = v3_1517448501_843 == v3_1517448501_1003;
   assign v3_1517448501_1014 = a_c1 & v3_1517448501_1013;
   assign v3_1517448501_1015 = ~v3_1517448501_1016;
   assign v3_1517448501_1016 = f15 & ~v3_1517448501_1014;
   assign v3_1517448501_1017 = v3_1517448501_1002 & v3_1517448501_1015;
   assign v3_1517448501_1018 = v3_1517448501_930 == v3_1517448501_1003;
   assign v3_1517448501_1019 = a_c1 & v3_1517448501_1018;
   assign v3_1517448501_1020 = ~v3_1517448501_1021;
   assign v3_1517448501_1021 = f16 & ~v3_1517448501_1019;
   assign v3_1517448501_1022 = v3_1517448501_1017 & v3_1517448501_1020;
   assign v3_1517448501_1023 = ~v3_1517448501_1013 & ~v3_1517448501_1018;
   assign v3_1517448501_1024 = a_c1 & v3_1517448501_1023;
   assign v3_1517448501_1025 = ~v3_1517448501_1026;
   assign v3_1517448501_1026 = f17 & ~v3_1517448501_1024;
   assign v3_1517448501_1027 = v3_1517448501_1022 & v3_1517448501_1025;
   assign v3_1517448501_1028 = v3_1517448501_1029 ? v3_1517448501_1037 : v3_1517448501_1036;
   assign v3_1517448501_1029 = v3_1517448501_979[31];
   assign v3_1517448501_1030 = v3_1517448501_111[31];
   assign v3_1517448501_1031 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1032 = ~v3_1517448501_979 + v3_1517448501_1031;
   assign v3_1517448501_1033 = ~v3_1517448501_111 + v3_1517448501_1031;
   assign v3_1517448501_1034 = v3_1517448501_1029 ? v3_1517448501_1032 : v3_1517448501_979;
   assign v3_1517448501_1035 = v3_1517448501_1030 ? v3_1517448501_1033 : v3_1517448501_111;
   assign v3_1517448501_1036 = v3_1517448501_1034 % v3_1517448501_1035;
   assign v3_1517448501_1037 = ~v3_1517448501_1036 + v3_1517448501_1031;
   assign v3_1517448501_1038 = v3_1517448501_1041 ? v3_1517448501_1048 : v3_1517448501_1047;
   assign v3_1517448501_1039 = v3_1517448501_1028[31];
   assign v3_1517448501_1040 = v3_1517448501_77[31];
   assign v3_1517448501_1041 = v3_1517448501_1039 ^ v3_1517448501_1040;
   assign v3_1517448501_1042 = 32'b00000000_00000000_00000000_00000001; 
   assign v3_1517448501_1043 = ~v3_1517448501_1028 + v3_1517448501_1042;
   assign v3_1517448501_1044 = ~v3_1517448501_77 + v3_1517448501_1042;
   assign v3_1517448501_1045 = v3_1517448501_1039 ? v3_1517448501_1043 : v3_1517448501_1028;
   assign v3_1517448501_1046 = v3_1517448501_1040 ? v3_1517448501_1044 : v3_1517448501_77;
   assign v3_1517448501_1047 = v3_1517448501_1045 / v3_1517448501_1046;
   assign v3_1517448501_1048 = ~v3_1517448501_1047 + v3_1517448501_1042;
   assign v3_1517448501_1049 = v3_1517448501_909 == v3_1517448501_1038;
   assign v3_1517448501_1050 = v3_1517448501_1018 & v3_1517448501_1049;
   assign v3_1517448501_1051 = a_c2 & v3_1517448501_1050;
   assign v3_1517448501_1052 = ~v3_1517448501_1053;
   assign v3_1517448501_1053 = f18 & ~v3_1517448501_1051;
   assign v3_1517448501_1054 = v3_1517448501_1027 & v3_1517448501_1052;
   assign v3_1517448501_1055 = a_c2 & ~v3_1517448501_1050;
   assign v3_1517448501_1056 = ~v3_1517448501_1057;
   assign v3_1517448501_1057 = f19 & ~v3_1517448501_1055;
   assign v3_1517448501_1058 = v3_1517448501_1054 & v3_1517448501_1056;
   assign v3_1517448501_1059 = v3_1517448501_52 == v3_1517448501_1038;
   assign v3_1517448501_1060 = v3_1517448501_1013 & v3_1517448501_1059;
   assign v3_1517448501_1061 = v3_1517448501_909 == v3_1517448501_983;
   assign v3_1517448501_1062 = v3_1517448501_1060 & v3_1517448501_1061;
   assign v3_1517448501_1063 = a_d1 & v3_1517448501_1062;
   assign v3_1517448501_1064 = ~v3_1517448501_1065;
   assign v3_1517448501_1065 = f20 & ~v3_1517448501_1063;
   assign v3_1517448501_1066 = v3_1517448501_1058 & v3_1517448501_1064;
   assign v3_1517448501_1067 = v3_1517448501_930 == v3_1517448501_1038;
   assign v3_1517448501_1068 = v3_1517448501_1013 & v3_1517448501_1067;
   assign v3_1517448501_1069 = v3_1517448501_52 == v3_1517448501_983;
   assign v3_1517448501_1070 = v3_1517448501_1068 & v3_1517448501_1069;
   assign v3_1517448501_1071 = a_d1 & v3_1517448501_1070;
   assign v3_1517448501_1072 = ~v3_1517448501_1073;
   assign v3_1517448501_1073 = f21 & ~v3_1517448501_1071;
   assign v3_1517448501_1074 = v3_1517448501_1066 & v3_1517448501_1072;
   assign v3_1517448501_1075 = ~v3_1517448501_1076;
   assign v3_1517448501_1076 = ~a_d1 & f22;
   assign v3_1517448501_1077 = v3_1517448501_1074 & v3_1517448501_1075;
   assign v3_1517448501_1078 = v3_1517448501_875 == v3_1517448501_1038;
   assign v3_1517448501_1079 = a_got2 & v3_1517448501_1078;
   assign v3_1517448501_1080 = ~v3_1517448501_1081;
   assign v3_1517448501_1081 = f23 & ~v3_1517448501_1079;
   assign v3_1517448501_1082 = v3_1517448501_1077 & v3_1517448501_1080;
   assign v3_1517448501_1083 = a_got2 & ~v3_1517448501_1078;
   assign v3_1517448501_1084 = ~v3_1517448501_1085;
   assign v3_1517448501_1085 = f24 & ~v3_1517448501_1083;
   assign v3_1517448501_1086 = v3_1517448501_1082 & v3_1517448501_1084;
   assign v3_1517448501_1087 = a_e1 & v3_1517448501_1013;
   assign v3_1517448501_1088 = ~v3_1517448501_1089;
   assign v3_1517448501_1089 = f25 & ~v3_1517448501_1087;
   assign v3_1517448501_1090 = v3_1517448501_1086 & v3_1517448501_1088;
   assign v3_1517448501_1091 = a_e1 & v3_1517448501_1018;
   assign v3_1517448501_1092 = ~v3_1517448501_1093;
   assign v3_1517448501_1093 = f26 & ~v3_1517448501_1091;
   assign v3_1517448501_1094 = v3_1517448501_1090 & v3_1517448501_1092;
   assign v3_1517448501_1095 = a_e1 & v3_1517448501_1023;
   assign v3_1517448501_1096 = ~v3_1517448501_1097;
   assign v3_1517448501_1097 = f27 & ~v3_1517448501_1095;
   assign v3_1517448501_1098 = v3_1517448501_1094 & v3_1517448501_1096;
   assign v3_1517448501_1099 = a_f1 & v3_1517448501_1050;
   assign v3_1517448501_1100 = ~v3_1517448501_1101;
   assign v3_1517448501_1101 = f28 & ~v3_1517448501_1099;
   assign v3_1517448501_1102 = v3_1517448501_1098 & v3_1517448501_1100;
   assign v3_1517448501_1103 = a_f1 & ~v3_1517448501_1050;
   assign v3_1517448501_1104 = ~v3_1517448501_1105;
   assign v3_1517448501_1105 = f29 & ~v3_1517448501_1103;
   assign v3_1517448501_1106 = v3_1517448501_1102 & v3_1517448501_1104;
   assign v3_1517448501_1107 = ~a_start_initiator_0 & ~a_start_responder_0;
   assign v3_1517448501_1108 = ~v3_1517448501_1109;
   assign v3_1517448501_1109 = f30 & ~v3_1517448501_1107;
   assign v3_1517448501_1110 = v3_1517448501_1106 & v3_1517448501_1108;
   assign v3_1517448501_1111 = ~a_start_initiator_0 & ~a_start_responder_1;
   assign v3_1517448501_1112 = ~v3_1517448501_1113;
   assign v3_1517448501_1113 = f31 & ~v3_1517448501_1111;
   assign v3_1517448501_1114 = v3_1517448501_1110 & v3_1517448501_1112;
   assign v3_1517448501_1115 = ~a_start_initiator_0 & ~a_q;
   assign v3_1517448501_1116 = ~v3_1517448501_1117;
   assign v3_1517448501_1117 = f32 & ~v3_1517448501_1115;
   assign v3_1517448501_1118 = v3_1517448501_1114 & v3_1517448501_1116;
   assign v3_1517448501_1119 = ~a_start_initiator_1 & ~a_start_responder_0;
   assign v3_1517448501_1120 = ~v3_1517448501_1121;
   assign v3_1517448501_1121 = f33 & ~v3_1517448501_1119;
   assign v3_1517448501_1122 = v3_1517448501_1118 & v3_1517448501_1120;
   assign v3_1517448501_1123 = ~a_start_initiator_1 & ~a_start_responder_1;
   assign v3_1517448501_1124 = ~v3_1517448501_1125;
   assign v3_1517448501_1125 = f34 & ~v3_1517448501_1123;
   assign v3_1517448501_1126 = v3_1517448501_1122 & v3_1517448501_1124;
   assign v3_1517448501_1127 = ~a_start_initiator_1 & ~a_q;
   assign v3_1517448501_1128 = ~v3_1517448501_1129;
   assign v3_1517448501_1129 = f35 & ~v3_1517448501_1127;
   assign v3_1517448501_1130 = v3_1517448501_1126 & v3_1517448501_1128;
   assign v3_1517448501_1131 = ~a_start_responder_0 & ~a_q;
   assign v3_1517448501_1132 = ~v3_1517448501_1133;
   assign v3_1517448501_1133 = f36 & ~v3_1517448501_1131;
   assign v3_1517448501_1134 = v3_1517448501_1130 & v3_1517448501_1132;
   assign v3_1517448501_1135 = ~a_start_responder_1 & ~a_q;
   assign v3_1517448501_1136 = ~v3_1517448501_1137;
   assign v3_1517448501_1137 = f37 & ~v3_1517448501_1135;
   assign v3_1517448501_1138 = v3_1517448501_1134 & v3_1517448501_1136;
   assign v3_1517448501_1139 = ~v3_1517448501_1140;
   assign v3_1517448501_1140 = ~v3_1517448501_1131 & f38;
   assign v3_1517448501_1141 = v3_1517448501_1138 & v3_1517448501_1139;
   assign v3_1517448501_1142 = ~v3_1517448501_1143;
   assign v3_1517448501_1143 = ~v3_1517448501_1135 & f39;
   assign v3_1517448501_1144 = v3_1517448501_1141 & v3_1517448501_1142;
   assign v3_1517448501_1145 = ~v3_1517448501_1146;
   assign v3_1517448501_1146 = ~v3_1517448501_1131 & f40;
   assign v3_1517448501_1147 = v3_1517448501_1144 & v3_1517448501_1145;
   assign v3_1517448501_1148 = ~v3_1517448501_1149;
   assign v3_1517448501_1149 = ~v3_1517448501_1135 & f41;
   assign v3_1517448501_1150 = v3_1517448501_1147 & v3_1517448501_1148;
   assign v3_1517448501_1151 = ~v3_1517448501_1152;
   assign v3_1517448501_1152 = ~v3_1517448501_1131 & f42;
   assign v3_1517448501_1153 = v3_1517448501_1150 & v3_1517448501_1151;
   assign v3_1517448501_1154 = ~v3_1517448501_1155;
   assign v3_1517448501_1155 = ~v3_1517448501_1135 & f43;
   assign v3_1517448501_1156 = v3_1517448501_1153 & v3_1517448501_1154;
   assign v3_1517448501_1157 = ~v3_1517448501_1158;
   assign v3_1517448501_1158 = ~v3_1517448501_1131 & f44;
   assign v3_1517448501_1159 = v3_1517448501_1156 & v3_1517448501_1157;
   assign v3_1517448501_1160 = ~v3_1517448501_1161;
   assign v3_1517448501_1161 = ~v3_1517448501_1135 & f45;
   assign v3_1517448501_1162 = v3_1517448501_1159 & v3_1517448501_1160;
   assign v3_1517448501_1163 = ~v3_1517448501_1164;
   assign v3_1517448501_1164 = ~v3_1517448501_1131 & f46;
   assign v3_1517448501_1165 = v3_1517448501_1162 & v3_1517448501_1163;
   assign v3_1517448501_1166 = ~v3_1517448501_1167;
   assign v3_1517448501_1167 = ~v3_1517448501_1135 & f47;
   assign v3_1517448501_1168 = v3_1517448501_1165 & v3_1517448501_1166;
   assign v3_1517448501_1169 = ~v3_1517448501_1170;
   assign v3_1517448501_1170 = ~v3_1517448501_1131 & f48;
   assign v3_1517448501_1171 = v3_1517448501_1168 & v3_1517448501_1169;
   assign v3_1517448501_1172 = ~v3_1517448501_1173;
   assign v3_1517448501_1173 = ~v3_1517448501_1135 & f49;
   assign v3_1517448501_1174 = v3_1517448501_1171 & v3_1517448501_1172;
   assign v3_1517448501_1175 = ~v3_1517448501_1176;
   assign v3_1517448501_1176 = ~v3_1517448501_1131 & f50;
   assign v3_1517448501_1177 = v3_1517448501_1174 & v3_1517448501_1175;
   assign v3_1517448501_1178 = ~v3_1517448501_1179;
   assign v3_1517448501_1179 = ~v3_1517448501_1135 & f51;
   assign v3_1517448501_1180 = v3_1517448501_1177 & v3_1517448501_1178;
   assign v3_1517448501_1181 = ~v3_1517448501_1182;
   assign v3_1517448501_1182 = ~v3_1517448501_1131 & f52;
   assign v3_1517448501_1183 = v3_1517448501_1180 & v3_1517448501_1181;
   assign v3_1517448501_1184 = ~v3_1517448501_1185;
   assign v3_1517448501_1185 = ~v3_1517448501_1135 & f53;
   assign v3_1517448501_1186 = v3_1517448501_1183 & v3_1517448501_1184;
   assign v3_1517448501_1187 = ~v3_1517448501_1188;
   assign v3_1517448501_1188 = ~v3_1517448501_1131 & f54;
   assign v3_1517448501_1189 = v3_1517448501_1186 & v3_1517448501_1187;
   assign v3_1517448501_1190 = ~v3_1517448501_1191;
   assign v3_1517448501_1191 = ~v3_1517448501_1135 & f55;
   assign v3_1517448501_1192 = v3_1517448501_1189 & v3_1517448501_1190;
   assign v3_1517448501_1193 = ~v3_1517448501_1194;
   assign v3_1517448501_1194 = ~v3_1517448501_1131 & f56;
   assign v3_1517448501_1195 = v3_1517448501_1192 & v3_1517448501_1193;
   assign v3_1517448501_1196 = ~v3_1517448501_1197;
   assign v3_1517448501_1197 = ~v3_1517448501_1135 & f57;
   assign v3_1517448501_1198 = v3_1517448501_1195 & v3_1517448501_1196;
   assign v3_1517448501_1199 = ~v3_1517448501_1200;
   assign v3_1517448501_1200 = ~v3_1517448501_1131 & f58;
   assign v3_1517448501_1201 = v3_1517448501_1198 & v3_1517448501_1199;
   assign v3_1517448501_1202 = ~v3_1517448501_1203;
   assign v3_1517448501_1203 = ~v3_1517448501_1135 & f59;
   assign v3_1517448501_1204 = v3_1517448501_1201 & v3_1517448501_1202;
   assign v3_1517448501_1205 = ~a_start_responder_0 & ~a_q;
   assign v3_1517448501_1206 = v3_1517448501_409 == v_kNa;
   assign v3_1517448501_1207 = v3_1517448501_1205 & v3_1517448501_1206;
   assign v3_1517448501_1208 = ~v3_1517448501_1209;
   assign v3_1517448501_1209 = f60 & ~v3_1517448501_1207;
   assign v3_1517448501_1210 = v3_1517448501_1204 & v3_1517448501_1208;
   assign v3_1517448501_1211 = ~a_start_responder_1 & ~a_q;
   assign v3_1517448501_1212 = v3_1517448501_1211 & v3_1517448501_1206;
   assign v3_1517448501_1213 = ~v3_1517448501_1214;
   assign v3_1517448501_1214 = f61 & ~v3_1517448501_1212;
   assign v3_1517448501_1215 = v3_1517448501_1210 & v3_1517448501_1213;
   assign v3_1517448501_1216 = ~v3_1517448501_1217;
   assign v3_1517448501_1217 = ~v3_1517448501_1207 & f62;
   assign v3_1517448501_1218 = v3_1517448501_1215 & v3_1517448501_1216;
   assign v3_1517448501_1219 = ~v3_1517448501_1220;
   assign v3_1517448501_1220 = ~v3_1517448501_1212 & f63;
   assign v3_1517448501_1221 = v3_1517448501_1218 & v3_1517448501_1219;
   assign v3_1517448501_1222 = ~v3_1517448501_1223;
   assign v3_1517448501_1223 = ~v3_1517448501_1207 & f64;
   assign v3_1517448501_1224 = v3_1517448501_1221 & v3_1517448501_1222;
   assign v3_1517448501_1225 = ~v3_1517448501_1226;
   assign v3_1517448501_1226 = ~v3_1517448501_1212 & f65;
   assign v3_1517448501_1227 = v3_1517448501_1224 & v3_1517448501_1225;
   assign v3_1517448501_1228 = ~a_start_responder_0 & ~a_q;
   assign v3_1517448501_1229 = 8'b00000000; 
   assign v3_1517448501_1230 = v3_1517448501_1229 == v_k_Na_A__B;
   assign v3_1517448501_1231 = ~v3_1517448501_1232;
   assign v3_1517448501_1232 = ~v3_1517448501_1206 & v3_1517448501_1230;
   assign v3_1517448501_1233 = v3_1517448501_1228 & v3_1517448501_1231;
   assign v3_1517448501_1234 = ~v3_1517448501_1235;
   assign v3_1517448501_1235 = f66 & ~v3_1517448501_1233;
   assign v3_1517448501_1236 = v3_1517448501_1227 & v3_1517448501_1234;
   assign v3_1517448501_1237 = ~a_start_responder_1 & ~a_q;
   assign v3_1517448501_1238 = v3_1517448501_1237 & v3_1517448501_1231;
   assign v3_1517448501_1239 = ~v3_1517448501_1240;
   assign v3_1517448501_1240 = f67 & ~v3_1517448501_1238;
   assign v3_1517448501_1241 = v3_1517448501_1236 & v3_1517448501_1239;
   assign v3_1517448501_1242 = ~v3_1517448501_1243;
   assign v3_1517448501_1243 = ~v3_1517448501_1207 & f68;
   assign v3_1517448501_1244 = v3_1517448501_1241 & v3_1517448501_1242;
   assign v3_1517448501_1245 = ~v3_1517448501_1246;
   assign v3_1517448501_1246 = ~v3_1517448501_1212 & f69;
   assign v3_1517448501_1247 = v3_1517448501_1244 & v3_1517448501_1245;
   assign v3_1517448501_1248 = ~v3_1517448501_1249;
   assign v3_1517448501_1249 = ~v3_1517448501_1207 & f70;
   assign v3_1517448501_1250 = v3_1517448501_1247 & v3_1517448501_1248;
   assign v3_1517448501_1251 = ~v3_1517448501_1252;
   assign v3_1517448501_1252 = ~v3_1517448501_1212 & f71;
   assign v3_1517448501_1253 = v3_1517448501_1250 & v3_1517448501_1251;
   assign v3_1517448501_1254 = ~a_start_responder_0 & ~a_q;
   assign v3_1517448501_1255 = v3_1517448501_409 == v_kNb;
   assign v3_1517448501_1256 = v3_1517448501_1254 & v3_1517448501_1255;
   assign v3_1517448501_1257 = ~v3_1517448501_1258;
   assign v3_1517448501_1258 = f72 & ~v3_1517448501_1256;
   assign v3_1517448501_1259 = v3_1517448501_1253 & v3_1517448501_1257;
   assign v3_1517448501_1260 = ~a_start_responder_1 & ~a_q;
   assign v3_1517448501_1261 = v3_1517448501_1260 & v3_1517448501_1255;
   assign v3_1517448501_1262 = ~v3_1517448501_1263;
   assign v3_1517448501_1263 = f73 & ~v3_1517448501_1261;
   assign v3_1517448501_1264 = v3_1517448501_1259 & v3_1517448501_1262;
   assign v3_1517448501_1265 = ~v3_1517448501_1266;
   assign v3_1517448501_1266 = ~v3_1517448501_1256 & f74;
   assign v3_1517448501_1267 = v3_1517448501_1264 & v3_1517448501_1265;
   assign v3_1517448501_1268 = ~v3_1517448501_1269;
   assign v3_1517448501_1269 = ~v3_1517448501_1261 & f75;
   assign v3_1517448501_1270 = v3_1517448501_1267 & v3_1517448501_1268;
   assign v3_1517448501_1271 = ~v3_1517448501_1272;
   assign v3_1517448501_1272 = ~v3_1517448501_1256 & f76;
   assign v3_1517448501_1273 = v3_1517448501_1270 & v3_1517448501_1271;
   assign v3_1517448501_1274 = ~v3_1517448501_1275;
   assign v3_1517448501_1275 = ~v3_1517448501_1261 & f77;
   assign v3_1517448501_1276 = v3_1517448501_1273 & v3_1517448501_1274;
   assign v3_1517448501_1277 = a_wait_resp_initiator_0 & a_send_reply_responder_0;
   assign v3_1517448501_1278 = ~v3_1517448501_1279;
   assign v3_1517448501_1279 = f78 & ~v3_1517448501_1277;
   assign v3_1517448501_1280 = v3_1517448501_1276 & v3_1517448501_1278;
   assign v3_1517448501_1281 = a_wait_resp_initiator_1 & a_send_reply_responder_0;
   assign v3_1517448501_1282 = ~v3_1517448501_1283;
   assign v3_1517448501_1283 = f79 & ~v3_1517448501_1281;
   assign v3_1517448501_1284 = v3_1517448501_1280 & v3_1517448501_1282;
   assign v3_1517448501_1285 = a_send_reply_responder_0 & ~a_q;
   assign v3_1517448501_1286 = ~v3_1517448501_1287;
   assign v3_1517448501_1287 = f80 & ~v3_1517448501_1285;
   assign v3_1517448501_1288 = v3_1517448501_1284 & v3_1517448501_1286;
   assign v3_1517448501_1289 = a_wait_resp_initiator_0 & a_send_reply_responder_1;
   assign v3_1517448501_1290 = ~v3_1517448501_1291;
   assign v3_1517448501_1291 = f81 & ~v3_1517448501_1289;
   assign v3_1517448501_1292 = v3_1517448501_1288 & v3_1517448501_1290;
   assign v3_1517448501_1293 = a_wait_resp_initiator_1 & a_send_reply_responder_1;
   assign v3_1517448501_1294 = ~v3_1517448501_1295;
   assign v3_1517448501_1295 = f82 & ~v3_1517448501_1293;
   assign v3_1517448501_1296 = v3_1517448501_1292 & v3_1517448501_1294;
   assign v3_1517448501_1297 = a_send_reply_responder_1 & ~a_q;
   assign v3_1517448501_1298 = ~v3_1517448501_1299;
   assign v3_1517448501_1299 = f83 & ~v3_1517448501_1297;
   assign v3_1517448501_1300 = v3_1517448501_1296 & v3_1517448501_1298;
   assign v3_1517448501_1301 = a_wait_resp_initiator_0 & ~a_q;
   assign v3_1517448501_1302 = v3_1517448501_1301 & v3_1517448501_1206;
   assign v3_1517448501_1303 = ~v3_1517448501_1304;
   assign v3_1517448501_1304 = f84 & ~v3_1517448501_1302;
   assign v3_1517448501_1305 = v3_1517448501_1300 & v3_1517448501_1303;
   assign v3_1517448501_1306 = a_wait_resp_initiator_1 & ~a_q;
   assign v3_1517448501_1307 = v3_1517448501_1306 & v3_1517448501_1206;
   assign v3_1517448501_1308 = ~v3_1517448501_1309;
   assign v3_1517448501_1309 = f85 & ~v3_1517448501_1307;
   assign v3_1517448501_1310 = v3_1517448501_1305 & v3_1517448501_1308;
   assign v3_1517448501_1311 = a_wait_resp_initiator_0 & ~a_q;
   assign v3_1517448501_1312 = v3_1517448501_1206 & v3_1517448501_1255;
   assign v3_1517448501_1313 = v3_1517448501_409 == v_k_Na_Nb__A;
   assign v3_1517448501_1314 = ~v3_1517448501_1315;
   assign v3_1517448501_1315 = ~v3_1517448501_1312 & ~v3_1517448501_1313;
   assign v3_1517448501_1316 = v3_1517448501_1311 & v3_1517448501_1314;
   assign v3_1517448501_1317 = ~v3_1517448501_1318;
   assign v3_1517448501_1318 = f86 & ~v3_1517448501_1316;
   assign v3_1517448501_1319 = v3_1517448501_1310 & v3_1517448501_1317;
   assign v3_1517448501_1320 = a_wait_resp_initiator_1 & ~a_q;
   assign v3_1517448501_1321 = v3_1517448501_1320 & v3_1517448501_1314;
   assign v3_1517448501_1322 = ~v3_1517448501_1323;
   assign v3_1517448501_1323 = f87 & ~v3_1517448501_1321;
   assign v3_1517448501_1324 = v3_1517448501_1319 & v3_1517448501_1322;
   assign v3_1517448501_1325 = ~v3_1517448501_1326;
   assign v3_1517448501_1326 = ~v3_1517448501_1302 & f88;
   assign v3_1517448501_1327 = v3_1517448501_1324 & v3_1517448501_1325;
   assign v3_1517448501_1328 = ~v3_1517448501_1329;
   assign v3_1517448501_1329 = ~v3_1517448501_1307 & f89;
   assign v3_1517448501_1330 = v3_1517448501_1327 & v3_1517448501_1328;
   assign v3_1517448501_1331 = a_commited_initiator_0 & a_wait_resp_responder_0;
   assign v3_1517448501_1332 = ~v3_1517448501_1333;
   assign v3_1517448501_1333 = f90 & ~v3_1517448501_1331;
   assign v3_1517448501_1334 = v3_1517448501_1330 & v3_1517448501_1332;
   assign v3_1517448501_1335 = a_commited_initiator_0 & a_wait_resp_responder_1;
   assign v3_1517448501_1336 = ~v3_1517448501_1337;
   assign v3_1517448501_1337 = f91 & ~v3_1517448501_1335;
   assign v3_1517448501_1338 = v3_1517448501_1334 & v3_1517448501_1336;
   assign v3_1517448501_1339 = a_commited_initiator_0 & ~a_q;
   assign v3_1517448501_1340 = ~v3_1517448501_1341;
   assign v3_1517448501_1341 = f92 & ~v3_1517448501_1339;
   assign v3_1517448501_1342 = v3_1517448501_1338 & v3_1517448501_1340;
   assign v3_1517448501_1343 = a_commited_initiator_1 & a_wait_resp_responder_0;
   assign v3_1517448501_1344 = ~v3_1517448501_1345;
   assign v3_1517448501_1345 = f93 & ~v3_1517448501_1343;
   assign v3_1517448501_1346 = v3_1517448501_1342 & v3_1517448501_1344;
   assign v3_1517448501_1347 = a_commited_initiator_1 & a_wait_resp_responder_1;
   assign v3_1517448501_1348 = ~v3_1517448501_1349;
   assign v3_1517448501_1349 = f94 & ~v3_1517448501_1347;
   assign v3_1517448501_1350 = v3_1517448501_1346 & v3_1517448501_1348;
   assign v3_1517448501_1351 = a_commited_initiator_1 & ~a_q;
   assign v3_1517448501_1352 = ~v3_1517448501_1353;
   assign v3_1517448501_1353 = f95 & ~v3_1517448501_1351;
   assign v3_1517448501_1354 = v3_1517448501_1350 & v3_1517448501_1352;
   assign v3_1517448501_1355 = a_wait_resp_responder_0 & ~a_q;
   assign v3_1517448501_1356 = v3_1517448501_409 == v_k_Nb__B;
   assign v3_1517448501_1357 = ~v3_1517448501_1358;
   assign v3_1517448501_1358 = ~v3_1517448501_1255 & ~v3_1517448501_1356;
   assign v3_1517448501_1359 = v3_1517448501_1355 & v3_1517448501_1357;
   assign v3_1517448501_1360 = ~v3_1517448501_1361;
   assign v3_1517448501_1361 = f96 & ~v3_1517448501_1359;
   assign v3_1517448501_1362 = v3_1517448501_1354 & v3_1517448501_1360;
   assign v3_1517448501_1363 = a_wait_resp_responder_1 & ~a_q;
   assign v3_1517448501_1364 = v3_1517448501_1363 & v3_1517448501_1357;
   assign v3_1517448501_1365 = ~v3_1517448501_1366;
   assign v3_1517448501_1366 = f97 & ~v3_1517448501_1364;
   assign v3_1517448501_1367 = v3_1517448501_1362 & v3_1517448501_1365;
   assign v3_1517448501_1368 = ~v3_1517448501_1369;
   assign v3_1517448501_1369 = ~f00 & ~f01;
   assign v3_1517448501_1370 = ~v3_1517448501_1371;
   assign v3_1517448501_1371 = ~f02 & ~v3_1517448501_1368;
   assign v3_1517448501_1372 = ~v3_1517448501_1373;
   assign v3_1517448501_1373 = ~f03 & ~v3_1517448501_1370;
   assign v3_1517448501_1374 = ~v3_1517448501_1375;
   assign v3_1517448501_1375 = ~f04 & ~v3_1517448501_1372;
   assign v3_1517448501_1376 = ~v3_1517448501_1377;
   assign v3_1517448501_1377 = ~f05 & ~v3_1517448501_1374;
   assign v3_1517448501_1378 = ~v3_1517448501_1379;
   assign v3_1517448501_1379 = ~f06 & ~v3_1517448501_1376;
   assign v3_1517448501_1380 = ~v3_1517448501_1381;
   assign v3_1517448501_1381 = ~f07 & ~v3_1517448501_1378;
   assign v3_1517448501_1382 = ~v3_1517448501_1383;
   assign v3_1517448501_1383 = ~f08 & ~v3_1517448501_1380;
   assign v3_1517448501_1384 = ~v3_1517448501_1385;
   assign v3_1517448501_1385 = ~f09 & ~v3_1517448501_1382;
   assign v3_1517448501_1386 = ~v3_1517448501_1387;
   assign v3_1517448501_1387 = ~f10 & ~v3_1517448501_1384;
   assign v3_1517448501_1388 = ~v3_1517448501_1389;
   assign v3_1517448501_1389 = ~f11 & ~v3_1517448501_1386;
   assign v3_1517448501_1390 = ~v3_1517448501_1391;
   assign v3_1517448501_1391 = ~f12 & ~v3_1517448501_1388;
   assign v3_1517448501_1392 = ~v3_1517448501_1393;
   assign v3_1517448501_1393 = ~f13 & ~v3_1517448501_1390;
   assign v3_1517448501_1394 = ~v3_1517448501_1395;
   assign v3_1517448501_1395 = ~f14 & ~v3_1517448501_1392;
   assign v3_1517448501_1396 = ~v3_1517448501_1397;
   assign v3_1517448501_1397 = ~f15 & ~v3_1517448501_1394;
   assign v3_1517448501_1398 = ~v3_1517448501_1399;
   assign v3_1517448501_1399 = ~f16 & ~v3_1517448501_1396;
   assign v3_1517448501_1400 = ~v3_1517448501_1401;
   assign v3_1517448501_1401 = ~f17 & ~v3_1517448501_1398;
   assign v3_1517448501_1402 = ~v3_1517448501_1403;
   assign v3_1517448501_1403 = ~f18 & ~v3_1517448501_1400;
   assign v3_1517448501_1404 = ~v3_1517448501_1405;
   assign v3_1517448501_1405 = ~f19 & ~v3_1517448501_1402;
   assign v3_1517448501_1406 = ~v3_1517448501_1407;
   assign v3_1517448501_1407 = ~f20 & ~v3_1517448501_1404;
   assign v3_1517448501_1408 = ~v3_1517448501_1409;
   assign v3_1517448501_1409 = ~f21 & ~v3_1517448501_1406;
   assign v3_1517448501_1410 = ~v3_1517448501_1411;
   assign v3_1517448501_1411 = ~f22 & ~v3_1517448501_1408;
   assign v3_1517448501_1412 = ~v3_1517448501_1413;
   assign v3_1517448501_1413 = ~f23 & ~v3_1517448501_1410;
   assign v3_1517448501_1414 = ~v3_1517448501_1415;
   assign v3_1517448501_1415 = ~f24 & ~v3_1517448501_1412;
   assign v3_1517448501_1416 = ~v3_1517448501_1417;
   assign v3_1517448501_1417 = ~f25 & ~v3_1517448501_1414;
   assign v3_1517448501_1418 = ~v3_1517448501_1419;
   assign v3_1517448501_1419 = ~f26 & ~v3_1517448501_1416;
   assign v3_1517448501_1420 = ~v3_1517448501_1421;
   assign v3_1517448501_1421 = ~f27 & ~v3_1517448501_1418;
   assign v3_1517448501_1422 = ~v3_1517448501_1423;
   assign v3_1517448501_1423 = ~f28 & ~v3_1517448501_1420;
   assign v3_1517448501_1424 = ~v3_1517448501_1425;
   assign v3_1517448501_1425 = ~f29 & ~v3_1517448501_1422;
   assign v3_1517448501_1426 = ~v3_1517448501_1427;
   assign v3_1517448501_1427 = ~f30 & ~v3_1517448501_1424;
   assign v3_1517448501_1428 = ~v3_1517448501_1429;
   assign v3_1517448501_1429 = ~f31 & ~v3_1517448501_1426;
   assign v3_1517448501_1430 = ~v3_1517448501_1431;
   assign v3_1517448501_1431 = ~f32 & ~v3_1517448501_1428;
   assign v3_1517448501_1432 = ~v3_1517448501_1433;
   assign v3_1517448501_1433 = ~f33 & ~v3_1517448501_1430;
   assign v3_1517448501_1434 = ~v3_1517448501_1435;
   assign v3_1517448501_1435 = ~f34 & ~v3_1517448501_1432;
   assign v3_1517448501_1436 = ~v3_1517448501_1437;
   assign v3_1517448501_1437 = ~f35 & ~v3_1517448501_1434;
   assign v3_1517448501_1438 = ~v3_1517448501_1439;
   assign v3_1517448501_1439 = ~f36 & ~v3_1517448501_1436;
   assign v3_1517448501_1440 = ~v3_1517448501_1441;
   assign v3_1517448501_1441 = ~f37 & ~v3_1517448501_1438;
   assign v3_1517448501_1442 = ~v3_1517448501_1443;
   assign v3_1517448501_1443 = ~f38 & ~v3_1517448501_1440;
   assign v3_1517448501_1444 = ~v3_1517448501_1445;
   assign v3_1517448501_1445 = ~f39 & ~v3_1517448501_1442;
   assign v3_1517448501_1446 = ~v3_1517448501_1447;
   assign v3_1517448501_1447 = ~f40 & ~v3_1517448501_1444;
   assign v3_1517448501_1448 = ~v3_1517448501_1449;
   assign v3_1517448501_1449 = ~f41 & ~v3_1517448501_1446;
   assign v3_1517448501_1450 = ~v3_1517448501_1451;
   assign v3_1517448501_1451 = ~f42 & ~v3_1517448501_1448;
   assign v3_1517448501_1452 = ~v3_1517448501_1453;
   assign v3_1517448501_1453 = ~f43 & ~v3_1517448501_1450;
   assign v3_1517448501_1454 = ~v3_1517448501_1455;
   assign v3_1517448501_1455 = ~f44 & ~v3_1517448501_1452;
   assign v3_1517448501_1456 = ~v3_1517448501_1457;
   assign v3_1517448501_1457 = ~f45 & ~v3_1517448501_1454;
   assign v3_1517448501_1458 = ~v3_1517448501_1459;
   assign v3_1517448501_1459 = ~f46 & ~v3_1517448501_1456;
   assign v3_1517448501_1460 = ~v3_1517448501_1461;
   assign v3_1517448501_1461 = ~f47 & ~v3_1517448501_1458;
   assign v3_1517448501_1462 = ~v3_1517448501_1463;
   assign v3_1517448501_1463 = ~f48 & ~v3_1517448501_1460;
   assign v3_1517448501_1464 = ~v3_1517448501_1465;
   assign v3_1517448501_1465 = ~f49 & ~v3_1517448501_1462;
   assign v3_1517448501_1466 = ~v3_1517448501_1467;
   assign v3_1517448501_1467 = ~f50 & ~v3_1517448501_1464;
   assign v3_1517448501_1468 = ~v3_1517448501_1469;
   assign v3_1517448501_1469 = ~f51 & ~v3_1517448501_1466;
   assign v3_1517448501_1470 = ~v3_1517448501_1471;
   assign v3_1517448501_1471 = ~f52 & ~v3_1517448501_1468;
   assign v3_1517448501_1472 = ~v3_1517448501_1473;
   assign v3_1517448501_1473 = ~f53 & ~v3_1517448501_1470;
   assign v3_1517448501_1474 = ~v3_1517448501_1475;
   assign v3_1517448501_1475 = ~f54 & ~v3_1517448501_1472;
   assign v3_1517448501_1476 = ~v3_1517448501_1477;
   assign v3_1517448501_1477 = ~f55 & ~v3_1517448501_1474;
   assign v3_1517448501_1478 = ~v3_1517448501_1479;
   assign v3_1517448501_1479 = ~f56 & ~v3_1517448501_1476;
   assign v3_1517448501_1480 = ~v3_1517448501_1481;
   assign v3_1517448501_1481 = ~f57 & ~v3_1517448501_1478;
   assign v3_1517448501_1482 = ~v3_1517448501_1483;
   assign v3_1517448501_1483 = ~f58 & ~v3_1517448501_1480;
   assign v3_1517448501_1484 = ~v3_1517448501_1485;
   assign v3_1517448501_1485 = ~f59 & ~v3_1517448501_1482;
   assign v3_1517448501_1486 = ~v3_1517448501_1487;
   assign v3_1517448501_1487 = ~f60 & ~v3_1517448501_1484;
   assign v3_1517448501_1488 = ~v3_1517448501_1489;
   assign v3_1517448501_1489 = ~f61 & ~v3_1517448501_1486;
   assign v3_1517448501_1490 = ~v3_1517448501_1491;
   assign v3_1517448501_1491 = ~f62 & ~v3_1517448501_1488;
   assign v3_1517448501_1492 = ~v3_1517448501_1493;
   assign v3_1517448501_1493 = ~f63 & ~v3_1517448501_1490;
   assign v3_1517448501_1494 = ~v3_1517448501_1495;
   assign v3_1517448501_1495 = ~f64 & ~v3_1517448501_1492;
   assign v3_1517448501_1496 = ~v3_1517448501_1497;
   assign v3_1517448501_1497 = ~f65 & ~v3_1517448501_1494;
   assign v3_1517448501_1498 = ~v3_1517448501_1499;
   assign v3_1517448501_1499 = ~f66 & ~v3_1517448501_1496;
   assign v3_1517448501_1500 = ~v3_1517448501_1501;
   assign v3_1517448501_1501 = ~f67 & ~v3_1517448501_1498;
   assign v3_1517448501_1502 = ~v3_1517448501_1503;
   assign v3_1517448501_1503 = ~f68 & ~v3_1517448501_1500;
   assign v3_1517448501_1504 = ~v3_1517448501_1505;
   assign v3_1517448501_1505 = ~f69 & ~v3_1517448501_1502;
   assign v3_1517448501_1506 = ~v3_1517448501_1507;
   assign v3_1517448501_1507 = ~f70 & ~v3_1517448501_1504;
   assign v3_1517448501_1508 = ~v3_1517448501_1509;
   assign v3_1517448501_1509 = ~f71 & ~v3_1517448501_1506;
   assign v3_1517448501_1510 = ~v3_1517448501_1511;
   assign v3_1517448501_1511 = ~f72 & ~v3_1517448501_1508;
   assign v3_1517448501_1512 = ~v3_1517448501_1513;
   assign v3_1517448501_1513 = ~f73 & ~v3_1517448501_1510;
   assign v3_1517448501_1514 = ~v3_1517448501_1515;
   assign v3_1517448501_1515 = ~f74 & ~v3_1517448501_1512;
   assign v3_1517448501_1516 = ~v3_1517448501_1517;
   assign v3_1517448501_1517 = ~f75 & ~v3_1517448501_1514;
   assign v3_1517448501_1518 = ~v3_1517448501_1519;
   assign v3_1517448501_1519 = ~f76 & ~v3_1517448501_1516;
   assign v3_1517448501_1520 = ~v3_1517448501_1521;
   assign v3_1517448501_1521 = ~f77 & ~v3_1517448501_1518;
   assign v3_1517448501_1522 = ~v3_1517448501_1523;
   assign v3_1517448501_1523 = ~f78 & ~v3_1517448501_1520;
   assign v3_1517448501_1524 = ~v3_1517448501_1525;
   assign v3_1517448501_1525 = ~f79 & ~v3_1517448501_1522;
   assign v3_1517448501_1526 = ~v3_1517448501_1527;
   assign v3_1517448501_1527 = ~f80 & ~v3_1517448501_1524;
   assign v3_1517448501_1528 = ~v3_1517448501_1529;
   assign v3_1517448501_1529 = ~f81 & ~v3_1517448501_1526;
   assign v3_1517448501_1530 = ~v3_1517448501_1531;
   assign v3_1517448501_1531 = ~f82 & ~v3_1517448501_1528;
   assign v3_1517448501_1532 = ~v3_1517448501_1533;
   assign v3_1517448501_1533 = ~f83 & ~v3_1517448501_1530;
   assign v3_1517448501_1534 = ~v3_1517448501_1535;
   assign v3_1517448501_1535 = ~f84 & ~v3_1517448501_1532;
   assign v3_1517448501_1536 = ~v3_1517448501_1537;
   assign v3_1517448501_1537 = ~f85 & ~v3_1517448501_1534;
   assign v3_1517448501_1538 = ~v3_1517448501_1539;
   assign v3_1517448501_1539 = ~f86 & ~v3_1517448501_1536;
   assign v3_1517448501_1540 = ~v3_1517448501_1541;
   assign v3_1517448501_1541 = ~f87 & ~v3_1517448501_1538;
   assign v3_1517448501_1542 = ~v3_1517448501_1543;
   assign v3_1517448501_1543 = ~f88 & ~v3_1517448501_1540;
   assign v3_1517448501_1544 = ~v3_1517448501_1545;
   assign v3_1517448501_1545 = ~f89 & ~v3_1517448501_1542;
   assign v3_1517448501_1546 = ~v3_1517448501_1547;
   assign v3_1517448501_1547 = ~f90 & ~v3_1517448501_1544;
   assign v3_1517448501_1548 = ~v3_1517448501_1549;
   assign v3_1517448501_1549 = ~f91 & ~v3_1517448501_1546;
   assign v3_1517448501_1550 = ~v3_1517448501_1551;
   assign v3_1517448501_1551 = ~f92 & ~v3_1517448501_1548;
   assign v3_1517448501_1552 = ~v3_1517448501_1553;
   assign v3_1517448501_1553 = ~f93 & ~v3_1517448501_1550;
   assign v3_1517448501_1554 = ~v3_1517448501_1555;
   assign v3_1517448501_1555 = ~f94 & ~v3_1517448501_1552;
   assign v3_1517448501_1556 = ~v3_1517448501_1557;
   assign v3_1517448501_1557 = ~f95 & ~v3_1517448501_1554;
   assign v3_1517448501_1558 = ~v3_1517448501_1559;
   assign v3_1517448501_1559 = ~f96 & ~v3_1517448501_1556;
   assign v3_1517448501_1560 = ~v3_1517448501_1561;
   assign v3_1517448501_1561 = ~f97 & ~v3_1517448501_1558;
   assign v3_1517448501_1562 = v3_1517448501_1367 & v3_1517448501_1560;
   assign v3_1517448501_1563 = f00 & f01;
   assign v3_1517448501_1564 = f02 & v3_1517448501_1368;
   assign v3_1517448501_1565 = ~v3_1517448501_1566;
   assign v3_1517448501_1566 = ~v3_1517448501_1563 & ~v3_1517448501_1564;
   assign v3_1517448501_1567 = f03 & v3_1517448501_1370;
   assign v3_1517448501_1568 = ~v3_1517448501_1569;
   assign v3_1517448501_1569 = ~v3_1517448501_1565 & ~v3_1517448501_1567;
   assign v3_1517448501_1570 = f04 & v3_1517448501_1372;
   assign v3_1517448501_1571 = ~v3_1517448501_1572;
   assign v3_1517448501_1572 = ~v3_1517448501_1568 & ~v3_1517448501_1570;
   assign v3_1517448501_1573 = f05 & v3_1517448501_1374;
   assign v3_1517448501_1574 = ~v3_1517448501_1575;
   assign v3_1517448501_1575 = ~v3_1517448501_1571 & ~v3_1517448501_1573;
   assign v3_1517448501_1576 = f06 & v3_1517448501_1376;
   assign v3_1517448501_1577 = ~v3_1517448501_1578;
   assign v3_1517448501_1578 = ~v3_1517448501_1574 & ~v3_1517448501_1576;
   assign v3_1517448501_1579 = f07 & v3_1517448501_1378;
   assign v3_1517448501_1580 = ~v3_1517448501_1581;
   assign v3_1517448501_1581 = ~v3_1517448501_1577 & ~v3_1517448501_1579;
   assign v3_1517448501_1582 = f08 & v3_1517448501_1380;
   assign v3_1517448501_1583 = ~v3_1517448501_1584;
   assign v3_1517448501_1584 = ~v3_1517448501_1580 & ~v3_1517448501_1582;
   assign v3_1517448501_1585 = f09 & v3_1517448501_1382;
   assign v3_1517448501_1586 = ~v3_1517448501_1587;
   assign v3_1517448501_1587 = ~v3_1517448501_1583 & ~v3_1517448501_1585;
   assign v3_1517448501_1588 = f10 & v3_1517448501_1384;
   assign v3_1517448501_1589 = ~v3_1517448501_1590;
   assign v3_1517448501_1590 = ~v3_1517448501_1586 & ~v3_1517448501_1588;
   assign v3_1517448501_1591 = f11 & v3_1517448501_1386;
   assign v3_1517448501_1592 = ~v3_1517448501_1593;
   assign v3_1517448501_1593 = ~v3_1517448501_1589 & ~v3_1517448501_1591;
   assign v3_1517448501_1594 = f12 & v3_1517448501_1388;
   assign v3_1517448501_1595 = ~v3_1517448501_1596;
   assign v3_1517448501_1596 = ~v3_1517448501_1592 & ~v3_1517448501_1594;
   assign v3_1517448501_1597 = f13 & v3_1517448501_1390;
   assign v3_1517448501_1598 = ~v3_1517448501_1599;
   assign v3_1517448501_1599 = ~v3_1517448501_1595 & ~v3_1517448501_1597;
   assign v3_1517448501_1600 = f14 & v3_1517448501_1392;
   assign v3_1517448501_1601 = ~v3_1517448501_1602;
   assign v3_1517448501_1602 = ~v3_1517448501_1598 & ~v3_1517448501_1600;
   assign v3_1517448501_1603 = f15 & v3_1517448501_1394;
   assign v3_1517448501_1604 = ~v3_1517448501_1605;
   assign v3_1517448501_1605 = ~v3_1517448501_1601 & ~v3_1517448501_1603;
   assign v3_1517448501_1606 = f16 & v3_1517448501_1396;
   assign v3_1517448501_1607 = ~v3_1517448501_1608;
   assign v3_1517448501_1608 = ~v3_1517448501_1604 & ~v3_1517448501_1606;
   assign v3_1517448501_1609 = f17 & v3_1517448501_1398;
   assign v3_1517448501_1610 = ~v3_1517448501_1611;
   assign v3_1517448501_1611 = ~v3_1517448501_1607 & ~v3_1517448501_1609;
   assign v3_1517448501_1612 = f18 & v3_1517448501_1400;
   assign v3_1517448501_1613 = ~v3_1517448501_1614;
   assign v3_1517448501_1614 = ~v3_1517448501_1610 & ~v3_1517448501_1612;
   assign v3_1517448501_1615 = f19 & v3_1517448501_1402;
   assign v3_1517448501_1616 = ~v3_1517448501_1617;
   assign v3_1517448501_1617 = ~v3_1517448501_1613 & ~v3_1517448501_1615;
   assign v3_1517448501_1618 = f20 & v3_1517448501_1404;
   assign v3_1517448501_1619 = ~v3_1517448501_1620;
   assign v3_1517448501_1620 = ~v3_1517448501_1616 & ~v3_1517448501_1618;
   assign v3_1517448501_1621 = f21 & v3_1517448501_1406;
   assign v3_1517448501_1622 = ~v3_1517448501_1623;
   assign v3_1517448501_1623 = ~v3_1517448501_1619 & ~v3_1517448501_1621;
   assign v3_1517448501_1624 = f22 & v3_1517448501_1408;
   assign v3_1517448501_1625 = ~v3_1517448501_1626;
   assign v3_1517448501_1626 = ~v3_1517448501_1622 & ~v3_1517448501_1624;
   assign v3_1517448501_1627 = f23 & v3_1517448501_1410;
   assign v3_1517448501_1628 = ~v3_1517448501_1629;
   assign v3_1517448501_1629 = ~v3_1517448501_1625 & ~v3_1517448501_1627;
   assign v3_1517448501_1630 = f24 & v3_1517448501_1412;
   assign v3_1517448501_1631 = ~v3_1517448501_1632;
   assign v3_1517448501_1632 = ~v3_1517448501_1628 & ~v3_1517448501_1630;
   assign v3_1517448501_1633 = f25 & v3_1517448501_1414;
   assign v3_1517448501_1634 = ~v3_1517448501_1635;
   assign v3_1517448501_1635 = ~v3_1517448501_1631 & ~v3_1517448501_1633;
   assign v3_1517448501_1636 = f26 & v3_1517448501_1416;
   assign v3_1517448501_1637 = ~v3_1517448501_1638;
   assign v3_1517448501_1638 = ~v3_1517448501_1634 & ~v3_1517448501_1636;
   assign v3_1517448501_1639 = f27 & v3_1517448501_1418;
   assign v3_1517448501_1640 = ~v3_1517448501_1641;
   assign v3_1517448501_1641 = ~v3_1517448501_1637 & ~v3_1517448501_1639;
   assign v3_1517448501_1642 = f28 & v3_1517448501_1420;
   assign v3_1517448501_1643 = ~v3_1517448501_1644;
   assign v3_1517448501_1644 = ~v3_1517448501_1640 & ~v3_1517448501_1642;
   assign v3_1517448501_1645 = f29 & v3_1517448501_1422;
   assign v3_1517448501_1646 = ~v3_1517448501_1647;
   assign v3_1517448501_1647 = ~v3_1517448501_1643 & ~v3_1517448501_1645;
   assign v3_1517448501_1648 = f30 & v3_1517448501_1424;
   assign v3_1517448501_1649 = ~v3_1517448501_1650;
   assign v3_1517448501_1650 = ~v3_1517448501_1646 & ~v3_1517448501_1648;
   assign v3_1517448501_1651 = f31 & v3_1517448501_1426;
   assign v3_1517448501_1652 = ~v3_1517448501_1653;
   assign v3_1517448501_1653 = ~v3_1517448501_1649 & ~v3_1517448501_1651;
   assign v3_1517448501_1654 = f32 & v3_1517448501_1428;
   assign v3_1517448501_1655 = ~v3_1517448501_1656;
   assign v3_1517448501_1656 = ~v3_1517448501_1652 & ~v3_1517448501_1654;
   assign v3_1517448501_1657 = f33 & v3_1517448501_1430;
   assign v3_1517448501_1658 = ~v3_1517448501_1659;
   assign v3_1517448501_1659 = ~v3_1517448501_1655 & ~v3_1517448501_1657;
   assign v3_1517448501_1660 = f34 & v3_1517448501_1432;
   assign v3_1517448501_1661 = ~v3_1517448501_1662;
   assign v3_1517448501_1662 = ~v3_1517448501_1658 & ~v3_1517448501_1660;
   assign v3_1517448501_1663 = f35 & v3_1517448501_1434;
   assign v3_1517448501_1664 = ~v3_1517448501_1665;
   assign v3_1517448501_1665 = ~v3_1517448501_1661 & ~v3_1517448501_1663;
   assign v3_1517448501_1666 = f36 & v3_1517448501_1436;
   assign v3_1517448501_1667 = ~v3_1517448501_1668;
   assign v3_1517448501_1668 = ~v3_1517448501_1664 & ~v3_1517448501_1666;
   assign v3_1517448501_1669 = f37 & v3_1517448501_1438;
   assign v3_1517448501_1670 = ~v3_1517448501_1671;
   assign v3_1517448501_1671 = ~v3_1517448501_1667 & ~v3_1517448501_1669;
   assign v3_1517448501_1672 = f38 & v3_1517448501_1440;
   assign v3_1517448501_1673 = ~v3_1517448501_1674;
   assign v3_1517448501_1674 = ~v3_1517448501_1670 & ~v3_1517448501_1672;
   assign v3_1517448501_1675 = f39 & v3_1517448501_1442;
   assign v3_1517448501_1676 = ~v3_1517448501_1677;
   assign v3_1517448501_1677 = ~v3_1517448501_1673 & ~v3_1517448501_1675;
   assign v3_1517448501_1678 = f40 & v3_1517448501_1444;
   assign v3_1517448501_1679 = ~v3_1517448501_1680;
   assign v3_1517448501_1680 = ~v3_1517448501_1676 & ~v3_1517448501_1678;
   assign v3_1517448501_1681 = f41 & v3_1517448501_1446;
   assign v3_1517448501_1682 = ~v3_1517448501_1683;
   assign v3_1517448501_1683 = ~v3_1517448501_1679 & ~v3_1517448501_1681;
   assign v3_1517448501_1684 = f42 & v3_1517448501_1448;
   assign v3_1517448501_1685 = ~v3_1517448501_1686;
   assign v3_1517448501_1686 = ~v3_1517448501_1682 & ~v3_1517448501_1684;
   assign v3_1517448501_1687 = f43 & v3_1517448501_1450;
   assign v3_1517448501_1688 = ~v3_1517448501_1689;
   assign v3_1517448501_1689 = ~v3_1517448501_1685 & ~v3_1517448501_1687;
   assign v3_1517448501_1690 = f44 & v3_1517448501_1452;
   assign v3_1517448501_1691 = ~v3_1517448501_1692;
   assign v3_1517448501_1692 = ~v3_1517448501_1688 & ~v3_1517448501_1690;
   assign v3_1517448501_1693 = f45 & v3_1517448501_1454;
   assign v3_1517448501_1694 = ~v3_1517448501_1695;
   assign v3_1517448501_1695 = ~v3_1517448501_1691 & ~v3_1517448501_1693;
   assign v3_1517448501_1696 = f46 & v3_1517448501_1456;
   assign v3_1517448501_1697 = ~v3_1517448501_1698;
   assign v3_1517448501_1698 = ~v3_1517448501_1694 & ~v3_1517448501_1696;
   assign v3_1517448501_1699 = f47 & v3_1517448501_1458;
   assign v3_1517448501_1700 = ~v3_1517448501_1701;
   assign v3_1517448501_1701 = ~v3_1517448501_1697 & ~v3_1517448501_1699;
   assign v3_1517448501_1702 = f48 & v3_1517448501_1460;
   assign v3_1517448501_1703 = ~v3_1517448501_1704;
   assign v3_1517448501_1704 = ~v3_1517448501_1700 & ~v3_1517448501_1702;
   assign v3_1517448501_1705 = f49 & v3_1517448501_1462;
   assign v3_1517448501_1706 = ~v3_1517448501_1707;
   assign v3_1517448501_1707 = ~v3_1517448501_1703 & ~v3_1517448501_1705;
   assign v3_1517448501_1708 = f50 & v3_1517448501_1464;
   assign v3_1517448501_1709 = ~v3_1517448501_1710;
   assign v3_1517448501_1710 = ~v3_1517448501_1706 & ~v3_1517448501_1708;
   assign v3_1517448501_1711 = f51 & v3_1517448501_1466;
   assign v3_1517448501_1712 = ~v3_1517448501_1713;
   assign v3_1517448501_1713 = ~v3_1517448501_1709 & ~v3_1517448501_1711;
   assign v3_1517448501_1714 = f52 & v3_1517448501_1468;
   assign v3_1517448501_1715 = ~v3_1517448501_1716;
   assign v3_1517448501_1716 = ~v3_1517448501_1712 & ~v3_1517448501_1714;
   assign v3_1517448501_1717 = f53 & v3_1517448501_1470;
   assign v3_1517448501_1718 = ~v3_1517448501_1719;
   assign v3_1517448501_1719 = ~v3_1517448501_1715 & ~v3_1517448501_1717;
   assign v3_1517448501_1720 = f54 & v3_1517448501_1472;
   assign v3_1517448501_1721 = ~v3_1517448501_1722;
   assign v3_1517448501_1722 = ~v3_1517448501_1718 & ~v3_1517448501_1720;
   assign v3_1517448501_1723 = f55 & v3_1517448501_1474;
   assign v3_1517448501_1724 = ~v3_1517448501_1725;
   assign v3_1517448501_1725 = ~v3_1517448501_1721 & ~v3_1517448501_1723;
   assign v3_1517448501_1726 = f56 & v3_1517448501_1476;
   assign v3_1517448501_1727 = ~v3_1517448501_1728;
   assign v3_1517448501_1728 = ~v3_1517448501_1724 & ~v3_1517448501_1726;
   assign v3_1517448501_1729 = f57 & v3_1517448501_1478;
   assign v3_1517448501_1730 = ~v3_1517448501_1731;
   assign v3_1517448501_1731 = ~v3_1517448501_1727 & ~v3_1517448501_1729;
   assign v3_1517448501_1732 = f58 & v3_1517448501_1480;
   assign v3_1517448501_1733 = ~v3_1517448501_1734;
   assign v3_1517448501_1734 = ~v3_1517448501_1730 & ~v3_1517448501_1732;
   assign v3_1517448501_1735 = f59 & v3_1517448501_1482;
   assign v3_1517448501_1736 = ~v3_1517448501_1737;
   assign v3_1517448501_1737 = ~v3_1517448501_1733 & ~v3_1517448501_1735;
   assign v3_1517448501_1738 = f60 & v3_1517448501_1484;
   assign v3_1517448501_1739 = ~v3_1517448501_1740;
   assign v3_1517448501_1740 = ~v3_1517448501_1736 & ~v3_1517448501_1738;
   assign v3_1517448501_1741 = f61 & v3_1517448501_1486;
   assign v3_1517448501_1742 = ~v3_1517448501_1743;
   assign v3_1517448501_1743 = ~v3_1517448501_1739 & ~v3_1517448501_1741;
   assign v3_1517448501_1744 = f62 & v3_1517448501_1488;
   assign v3_1517448501_1745 = ~v3_1517448501_1746;
   assign v3_1517448501_1746 = ~v3_1517448501_1742 & ~v3_1517448501_1744;
   assign v3_1517448501_1747 = f63 & v3_1517448501_1490;
   assign v3_1517448501_1748 = ~v3_1517448501_1749;
   assign v3_1517448501_1749 = ~v3_1517448501_1745 & ~v3_1517448501_1747;
   assign v3_1517448501_1750 = f64 & v3_1517448501_1492;
   assign v3_1517448501_1751 = ~v3_1517448501_1752;
   assign v3_1517448501_1752 = ~v3_1517448501_1748 & ~v3_1517448501_1750;
   assign v3_1517448501_1753 = f65 & v3_1517448501_1494;
   assign v3_1517448501_1754 = ~v3_1517448501_1755;
   assign v3_1517448501_1755 = ~v3_1517448501_1751 & ~v3_1517448501_1753;
   assign v3_1517448501_1756 = f66 & v3_1517448501_1496;
   assign v3_1517448501_1757 = ~v3_1517448501_1758;
   assign v3_1517448501_1758 = ~v3_1517448501_1754 & ~v3_1517448501_1756;
   assign v3_1517448501_1759 = f67 & v3_1517448501_1498;
   assign v3_1517448501_1760 = ~v3_1517448501_1761;
   assign v3_1517448501_1761 = ~v3_1517448501_1757 & ~v3_1517448501_1759;
   assign v3_1517448501_1762 = f68 & v3_1517448501_1500;
   assign v3_1517448501_1763 = ~v3_1517448501_1764;
   assign v3_1517448501_1764 = ~v3_1517448501_1760 & ~v3_1517448501_1762;
   assign v3_1517448501_1765 = f69 & v3_1517448501_1502;
   assign v3_1517448501_1766 = ~v3_1517448501_1767;
   assign v3_1517448501_1767 = ~v3_1517448501_1763 & ~v3_1517448501_1765;
   assign v3_1517448501_1768 = f70 & v3_1517448501_1504;
   assign v3_1517448501_1769 = ~v3_1517448501_1770;
   assign v3_1517448501_1770 = ~v3_1517448501_1766 & ~v3_1517448501_1768;
   assign v3_1517448501_1771 = f71 & v3_1517448501_1506;
   assign v3_1517448501_1772 = ~v3_1517448501_1773;
   assign v3_1517448501_1773 = ~v3_1517448501_1769 & ~v3_1517448501_1771;
   assign v3_1517448501_1774 = f72 & v3_1517448501_1508;
   assign v3_1517448501_1775 = ~v3_1517448501_1776;
   assign v3_1517448501_1776 = ~v3_1517448501_1772 & ~v3_1517448501_1774;
   assign v3_1517448501_1777 = f73 & v3_1517448501_1510;
   assign v3_1517448501_1778 = ~v3_1517448501_1779;
   assign v3_1517448501_1779 = ~v3_1517448501_1775 & ~v3_1517448501_1777;
   assign v3_1517448501_1780 = f74 & v3_1517448501_1512;
   assign v3_1517448501_1781 = ~v3_1517448501_1782;
   assign v3_1517448501_1782 = ~v3_1517448501_1778 & ~v3_1517448501_1780;
   assign v3_1517448501_1783 = f75 & v3_1517448501_1514;
   assign v3_1517448501_1784 = ~v3_1517448501_1785;
   assign v3_1517448501_1785 = ~v3_1517448501_1781 & ~v3_1517448501_1783;
   assign v3_1517448501_1786 = f76 & v3_1517448501_1516;
   assign v3_1517448501_1787 = ~v3_1517448501_1788;
   assign v3_1517448501_1788 = ~v3_1517448501_1784 & ~v3_1517448501_1786;
   assign v3_1517448501_1789 = f77 & v3_1517448501_1518;
   assign v3_1517448501_1790 = ~v3_1517448501_1791;
   assign v3_1517448501_1791 = ~v3_1517448501_1787 & ~v3_1517448501_1789;
   assign v3_1517448501_1792 = f78 & v3_1517448501_1520;
   assign v3_1517448501_1793 = ~v3_1517448501_1794;
   assign v3_1517448501_1794 = ~v3_1517448501_1790 & ~v3_1517448501_1792;
   assign v3_1517448501_1795 = f79 & v3_1517448501_1522;
   assign v3_1517448501_1796 = ~v3_1517448501_1797;
   assign v3_1517448501_1797 = ~v3_1517448501_1793 & ~v3_1517448501_1795;
   assign v3_1517448501_1798 = f80 & v3_1517448501_1524;
   assign v3_1517448501_1799 = ~v3_1517448501_1800;
   assign v3_1517448501_1800 = ~v3_1517448501_1796 & ~v3_1517448501_1798;
   assign v3_1517448501_1801 = f81 & v3_1517448501_1526;
   assign v3_1517448501_1802 = ~v3_1517448501_1803;
   assign v3_1517448501_1803 = ~v3_1517448501_1799 & ~v3_1517448501_1801;
   assign v3_1517448501_1804 = f82 & v3_1517448501_1528;
   assign v3_1517448501_1805 = ~v3_1517448501_1806;
   assign v3_1517448501_1806 = ~v3_1517448501_1802 & ~v3_1517448501_1804;
   assign v3_1517448501_1807 = f83 & v3_1517448501_1530;
   assign v3_1517448501_1808 = ~v3_1517448501_1809;
   assign v3_1517448501_1809 = ~v3_1517448501_1805 & ~v3_1517448501_1807;
   assign v3_1517448501_1810 = f84 & v3_1517448501_1532;
   assign v3_1517448501_1811 = ~v3_1517448501_1812;
   assign v3_1517448501_1812 = ~v3_1517448501_1808 & ~v3_1517448501_1810;
   assign v3_1517448501_1813 = f85 & v3_1517448501_1534;
   assign v3_1517448501_1814 = ~v3_1517448501_1815;
   assign v3_1517448501_1815 = ~v3_1517448501_1811 & ~v3_1517448501_1813;
   assign v3_1517448501_1816 = f86 & v3_1517448501_1536;
   assign v3_1517448501_1817 = ~v3_1517448501_1818;
   assign v3_1517448501_1818 = ~v3_1517448501_1814 & ~v3_1517448501_1816;
   assign v3_1517448501_1819 = f87 & v3_1517448501_1538;
   assign v3_1517448501_1820 = ~v3_1517448501_1821;
   assign v3_1517448501_1821 = ~v3_1517448501_1817 & ~v3_1517448501_1819;
   assign v3_1517448501_1822 = f88 & v3_1517448501_1540;
   assign v3_1517448501_1823 = ~v3_1517448501_1824;
   assign v3_1517448501_1824 = ~v3_1517448501_1820 & ~v3_1517448501_1822;
   assign v3_1517448501_1825 = f89 & v3_1517448501_1542;
   assign v3_1517448501_1826 = ~v3_1517448501_1827;
   assign v3_1517448501_1827 = ~v3_1517448501_1823 & ~v3_1517448501_1825;
   assign v3_1517448501_1828 = f90 & v3_1517448501_1544;
   assign v3_1517448501_1829 = ~v3_1517448501_1830;
   assign v3_1517448501_1830 = ~v3_1517448501_1826 & ~v3_1517448501_1828;
   assign v3_1517448501_1831 = f91 & v3_1517448501_1546;
   assign v3_1517448501_1832 = ~v3_1517448501_1833;
   assign v3_1517448501_1833 = ~v3_1517448501_1829 & ~v3_1517448501_1831;
   assign v3_1517448501_1834 = f92 & v3_1517448501_1548;
   assign v3_1517448501_1835 = ~v3_1517448501_1836;
   assign v3_1517448501_1836 = ~v3_1517448501_1832 & ~v3_1517448501_1834;
   assign v3_1517448501_1837 = f93 & v3_1517448501_1550;
   assign v3_1517448501_1838 = ~v3_1517448501_1839;
   assign v3_1517448501_1839 = ~v3_1517448501_1835 & ~v3_1517448501_1837;
   assign v3_1517448501_1840 = f94 & v3_1517448501_1552;
   assign v3_1517448501_1841 = ~v3_1517448501_1842;
   assign v3_1517448501_1842 = ~v3_1517448501_1838 & ~v3_1517448501_1840;
   assign v3_1517448501_1843 = f95 & v3_1517448501_1554;
   assign v3_1517448501_1844 = ~v3_1517448501_1845;
   assign v3_1517448501_1845 = ~v3_1517448501_1841 & ~v3_1517448501_1843;
   assign v3_1517448501_1846 = f96 & v3_1517448501_1556;
   assign v3_1517448501_1847 = ~v3_1517448501_1848;
   assign v3_1517448501_1848 = ~v3_1517448501_1844 & ~v3_1517448501_1846;
   assign v3_1517448501_1849 = f97 & v3_1517448501_1558;
   assign v3_1517448501_1850 = ~v3_1517448501_1851;
   assign v3_1517448501_1851 = ~v3_1517448501_1847 & ~v3_1517448501_1849;
   assign v3_1517448501_1852 = v3_1517448501_1562 & ~v3_1517448501_1850;
   assign v3_1517448501_1853 = ~a_start_initiator_0 & a_wait_resp_initiator_0;
   assign v3_1517448501_1854 = ~v3_1517448501_1855;
   assign v3_1517448501_1855 = a_start_initiator_0 & ~a_wait_resp_initiator_0;
   assign v3_1517448501_1856 = a_got_resp_initiator_0 & v3_1517448501_1854;
   assign v3_1517448501_1857 = ~v3_1517448501_1858;
   assign v3_1517448501_1858 = ~v3_1517448501_1853 & ~v3_1517448501_1856;
   assign v3_1517448501_1859 = ~v3_1517448501_1860;
   assign v3_1517448501_1860 = ~a_got_resp_initiator_0 & ~v3_1517448501_1854;
   assign v3_1517448501_1861 = a_commited_initiator_0 & v3_1517448501_1859;
   assign v3_1517448501_1862 = ~v3_1517448501_1863;
   assign v3_1517448501_1863 = ~v3_1517448501_1857 & ~v3_1517448501_1861;
   assign v3_1517448501_1864 = ~v3_1517448501_1865;
   assign v3_1517448501_1865 = ~a_commited_initiator_0 & ~v3_1517448501_1859;
   assign v3_1517448501_1866 = a_finished_initiator_0 & v3_1517448501_1864;
   assign v3_1517448501_1867 = ~v3_1517448501_1868;
   assign v3_1517448501_1868 = ~v3_1517448501_1862 & ~v3_1517448501_1866;
   assign v3_1517448501_1869 = ~v3_1517448501_1870;
   assign v3_1517448501_1870 = ~a_finished_initiator_0 & ~v3_1517448501_1864;
   assign v3_1517448501_1871 = a_corrupted_initiator_0 & v3_1517448501_1869;
   assign v3_1517448501_1872 = ~v3_1517448501_1873;
   assign v3_1517448501_1873 = ~v3_1517448501_1867 & ~v3_1517448501_1871;
   assign v3_1517448501_1874 = ~v3_1517448501_1875;
   assign v3_1517448501_1875 = ~a_corrupted_initiator_0 & ~v3_1517448501_1869;
   assign v3_1517448501_1876 = ~v3_1517448501_1872 & v3_1517448501_1874;
   assign v3_1517448501_1877 = ~a_start_initiator_1 & a_wait_resp_initiator_1;
   assign v3_1517448501_1878 = ~v3_1517448501_1879;
   assign v3_1517448501_1879 = a_start_initiator_1 & ~a_wait_resp_initiator_1;
   assign v3_1517448501_1880 = a_got_resp_initiator_1 & v3_1517448501_1878;
   assign v3_1517448501_1881 = ~v3_1517448501_1882;
   assign v3_1517448501_1882 = ~v3_1517448501_1877 & ~v3_1517448501_1880;
   assign v3_1517448501_1883 = ~v3_1517448501_1884;
   assign v3_1517448501_1884 = ~a_got_resp_initiator_1 & ~v3_1517448501_1878;
   assign v3_1517448501_1885 = a_commited_initiator_1 & v3_1517448501_1883;
   assign v3_1517448501_1886 = ~v3_1517448501_1887;
   assign v3_1517448501_1887 = ~v3_1517448501_1881 & ~v3_1517448501_1885;
   assign v3_1517448501_1888 = ~v3_1517448501_1889;
   assign v3_1517448501_1889 = ~a_commited_initiator_1 & ~v3_1517448501_1883;
   assign v3_1517448501_1890 = a_finished_initiator_1 & v3_1517448501_1888;
   assign v3_1517448501_1891 = ~v3_1517448501_1892;
   assign v3_1517448501_1892 = ~v3_1517448501_1886 & ~v3_1517448501_1890;
   assign v3_1517448501_1893 = ~v3_1517448501_1894;
   assign v3_1517448501_1894 = ~a_finished_initiator_1 & ~v3_1517448501_1888;
   assign v3_1517448501_1895 = a_corrupted_initiator_1 & v3_1517448501_1893;
   assign v3_1517448501_1896 = ~v3_1517448501_1897;
   assign v3_1517448501_1897 = ~v3_1517448501_1891 & ~v3_1517448501_1895;
   assign v3_1517448501_1898 = v3_1517448501_1876 & ~v3_1517448501_1896;
   assign v3_1517448501_1899 = ~v3_1517448501_1900;
   assign v3_1517448501_1900 = ~a_corrupted_initiator_1 & ~v3_1517448501_1893;
   assign v3_1517448501_1901 = v3_1517448501_1898 & v3_1517448501_1899;
   assign v3_1517448501_1902 = ~a_start_responder_0 & a_got_msg_responder_0;
   assign v3_1517448501_1903 = ~v3_1517448501_1904;
   assign v3_1517448501_1904 = a_start_responder_0 & ~a_got_msg_responder_0;
   assign v3_1517448501_1905 = a_send_reply_responder_0 & v3_1517448501_1903;
   assign v3_1517448501_1906 = ~v3_1517448501_1907;
   assign v3_1517448501_1907 = ~v3_1517448501_1902 & ~v3_1517448501_1905;
   assign v3_1517448501_1908 = ~v3_1517448501_1909;
   assign v3_1517448501_1909 = ~a_send_reply_responder_0 & ~v3_1517448501_1903;
   assign v3_1517448501_1910 = a_wait_resp_responder_0 & v3_1517448501_1908;
   assign v3_1517448501_1911 = ~v3_1517448501_1912;
   assign v3_1517448501_1912 = ~v3_1517448501_1906 & ~v3_1517448501_1910;
   assign v3_1517448501_1913 = ~v3_1517448501_1914;
   assign v3_1517448501_1914 = ~a_wait_resp_responder_0 & ~v3_1517448501_1908;
   assign v3_1517448501_1915 = a_got_resp_responder_0 & v3_1517448501_1913;
   assign v3_1517448501_1916 = ~v3_1517448501_1917;
   assign v3_1517448501_1917 = ~v3_1517448501_1911 & ~v3_1517448501_1915;
   assign v3_1517448501_1918 = ~v3_1517448501_1919;
   assign v3_1517448501_1919 = ~a_got_resp_responder_0 & ~v3_1517448501_1913;
   assign v3_1517448501_1920 = a_finished_responder_0 & v3_1517448501_1918;
   assign v3_1517448501_1921 = ~v3_1517448501_1922;
   assign v3_1517448501_1922 = ~v3_1517448501_1916 & ~v3_1517448501_1920;
   assign v3_1517448501_1923 = ~v3_1517448501_1924;
   assign v3_1517448501_1924 = ~a_finished_responder_0 & ~v3_1517448501_1918;
   assign v3_1517448501_1925 = a_corrupted_responder_0 & v3_1517448501_1923;
   assign v3_1517448501_1926 = ~v3_1517448501_1927;
   assign v3_1517448501_1927 = ~v3_1517448501_1921 & ~v3_1517448501_1925;
   assign v3_1517448501_1928 = v3_1517448501_1901 & ~v3_1517448501_1926;
   assign v3_1517448501_1929 = ~v3_1517448501_1930;
   assign v3_1517448501_1930 = ~a_corrupted_responder_0 & ~v3_1517448501_1923;
   assign v3_1517448501_1931 = v3_1517448501_1928 & v3_1517448501_1929;
   assign v3_1517448501_1932 = ~a_start_responder_1 & a_got_msg_responder_1;
   assign v3_1517448501_1933 = ~v3_1517448501_1934;
   assign v3_1517448501_1934 = a_start_responder_1 & ~a_got_msg_responder_1;
   assign v3_1517448501_1935 = a_send_reply_responder_1 & v3_1517448501_1933;
   assign v3_1517448501_1936 = ~v3_1517448501_1937;
   assign v3_1517448501_1937 = ~v3_1517448501_1932 & ~v3_1517448501_1935;
   assign v3_1517448501_1938 = ~v3_1517448501_1939;
   assign v3_1517448501_1939 = ~a_send_reply_responder_1 & ~v3_1517448501_1933;
   assign v3_1517448501_1940 = a_wait_resp_responder_1 & v3_1517448501_1938;
   assign v3_1517448501_1941 = ~v3_1517448501_1942;
   assign v3_1517448501_1942 = ~v3_1517448501_1936 & ~v3_1517448501_1940;
   assign v3_1517448501_1943 = ~v3_1517448501_1944;
   assign v3_1517448501_1944 = ~a_wait_resp_responder_1 & ~v3_1517448501_1938;
   assign v3_1517448501_1945 = a_got_resp_responder_1 & v3_1517448501_1943;
   assign v3_1517448501_1946 = ~v3_1517448501_1947;
   assign v3_1517448501_1947 = ~v3_1517448501_1941 & ~v3_1517448501_1945;
   assign v3_1517448501_1948 = ~v3_1517448501_1949;
   assign v3_1517448501_1949 = ~a_got_resp_responder_1 & ~v3_1517448501_1943;
   assign v3_1517448501_1950 = a_finished_responder_1 & v3_1517448501_1948;
   assign v3_1517448501_1951 = ~v3_1517448501_1952;
   assign v3_1517448501_1952 = ~v3_1517448501_1946 & ~v3_1517448501_1950;
   assign v3_1517448501_1953 = ~v3_1517448501_1954;
   assign v3_1517448501_1954 = ~a_finished_responder_1 & ~v3_1517448501_1948;
   assign v3_1517448501_1955 = a_corrupted_responder_1 & v3_1517448501_1953;
   assign v3_1517448501_1956 = ~v3_1517448501_1957;
   assign v3_1517448501_1957 = ~v3_1517448501_1951 & ~v3_1517448501_1955;
   assign v3_1517448501_1958 = v3_1517448501_1931 & ~v3_1517448501_1956;
   assign v3_1517448501_1959 = ~v3_1517448501_1960;
   assign v3_1517448501_1960 = ~a_corrupted_responder_1 & ~v3_1517448501_1953;
   assign v3_1517448501_1961 = v3_1517448501_1958 & v3_1517448501_1959;
   assign v3_1517448501_1962 = ~a_q & a_got3;
   assign v3_1517448501_1963 = ~v3_1517448501_1964;
   assign v3_1517448501_1964 = a_q & ~a_got3;
   assign v3_1517448501_1965 = a_c1 & v3_1517448501_1963;
   assign v3_1517448501_1966 = ~v3_1517448501_1967;
   assign v3_1517448501_1967 = ~v3_1517448501_1962 & ~v3_1517448501_1965;
   assign v3_1517448501_1968 = ~v3_1517448501_1969;
   assign v3_1517448501_1969 = ~a_c1 & ~v3_1517448501_1963;
   assign v3_1517448501_1970 = a_c2 & v3_1517448501_1968;
   assign v3_1517448501_1971 = ~v3_1517448501_1972;
   assign v3_1517448501_1972 = ~v3_1517448501_1966 & ~v3_1517448501_1970;
   assign v3_1517448501_1973 = ~v3_1517448501_1974;
   assign v3_1517448501_1974 = ~a_c2 & ~v3_1517448501_1968;
   assign v3_1517448501_1975 = a_d1 & v3_1517448501_1973;
   assign v3_1517448501_1976 = ~v3_1517448501_1977;
   assign v3_1517448501_1977 = ~v3_1517448501_1971 & ~v3_1517448501_1975;
   assign v3_1517448501_1978 = ~v3_1517448501_1979;
   assign v3_1517448501_1979 = ~a_d1 & ~v3_1517448501_1973;
   assign v3_1517448501_1980 = a_got2 & v3_1517448501_1978;
   assign v3_1517448501_1981 = ~v3_1517448501_1982;
   assign v3_1517448501_1982 = ~v3_1517448501_1976 & ~v3_1517448501_1980;
   assign v3_1517448501_1983 = ~v3_1517448501_1984;
   assign v3_1517448501_1984 = ~a_got2 & ~v3_1517448501_1978;
   assign v3_1517448501_1985 = a_e1 & v3_1517448501_1983;
   assign v3_1517448501_1986 = ~v3_1517448501_1987;
   assign v3_1517448501_1987 = ~v3_1517448501_1981 & ~v3_1517448501_1985;
   assign v3_1517448501_1988 = ~v3_1517448501_1989;
   assign v3_1517448501_1989 = ~a_e1 & ~v3_1517448501_1983;
   assign v3_1517448501_1990 = a_f1 & v3_1517448501_1988;
   assign v3_1517448501_1991 = ~v3_1517448501_1992;
   assign v3_1517448501_1992 = ~v3_1517448501_1986 & ~v3_1517448501_1990;
   assign v3_1517448501_1993 = v3_1517448501_1961 & ~v3_1517448501_1991;
   assign v3_1517448501_1994 = ~v3_1517448501_1995;
   assign v3_1517448501_1995 = ~a_f1 & ~v3_1517448501_1988;
   assign v3_1517448501_1996 = v3_1517448501_1993 & v3_1517448501_1994;
   assign v3_1517448501_1997 = v3_1517448501_1852 & v3_1517448501_1996;
   assign v3_1517448501_1998 = v3_1517448501_445 & v3_1517448501_457;
   assign v3_1517448501_1999 = ~v3_1517448501_2000;
   assign v3_1517448501_2000 = ~v3_1517448501_445 & ~v3_1517448501_457;
   assign v3_1517448501_2001 = v3_1517448501_470 & v3_1517448501_1999;
   assign v3_1517448501_2002 = ~v3_1517448501_2003;
   assign v3_1517448501_2003 = ~v3_1517448501_1998 & ~v3_1517448501_2001;
   assign v3_1517448501_2004 = ~v3_1517448501_2005;
   assign v3_1517448501_2005 = ~v3_1517448501_470 & ~v3_1517448501_1999;
   assign v3_1517448501_2006 = v3_1517448501_477 & v3_1517448501_2004;
   assign v3_1517448501_2007 = ~v3_1517448501_2008;
   assign v3_1517448501_2008 = ~v3_1517448501_2002 & ~v3_1517448501_2006;
   assign v3_1517448501_2009 = ~v3_1517448501_2010;
   assign v3_1517448501_2010 = ~v3_1517448501_477 & ~v3_1517448501_2004;
   assign v3_1517448501_2011 = v3_1517448501_483 & v3_1517448501_2009;
   assign v3_1517448501_2012 = ~v3_1517448501_2013;
   assign v3_1517448501_2013 = ~v3_1517448501_2007 & ~v3_1517448501_2011;
   assign v3_1517448501_2014 = ~v3_1517448501_2015;
   assign v3_1517448501_2015 = ~v3_1517448501_483 & ~v3_1517448501_2009;
   assign v3_1517448501_2016 = v3_1517448501_486 & v3_1517448501_2014;
   assign v3_1517448501_2017 = ~v3_1517448501_2018;
   assign v3_1517448501_2018 = ~v3_1517448501_2012 & ~v3_1517448501_2016;
   assign v3_1517448501_2019 = ~v3_1517448501_2020;
   assign v3_1517448501_2020 = ~v3_1517448501_486 & ~v3_1517448501_2014;
   assign v3_1517448501_2021 = ~v3_1517448501_2017 & v3_1517448501_2019;
   assign v3_1517448501_2022 = v3_1517448501_491 & v3_1517448501_503;
   assign v3_1517448501_2023 = ~v3_1517448501_2024;
   assign v3_1517448501_2024 = ~v3_1517448501_491 & ~v3_1517448501_503;
   assign v3_1517448501_2025 = v3_1517448501_516 & v3_1517448501_2023;
   assign v3_1517448501_2026 = ~v3_1517448501_2027;
   assign v3_1517448501_2027 = ~v3_1517448501_2022 & ~v3_1517448501_2025;
   assign v3_1517448501_2028 = ~v3_1517448501_2029;
   assign v3_1517448501_2029 = ~v3_1517448501_516 & ~v3_1517448501_2023;
   assign v3_1517448501_2030 = v3_1517448501_523 & v3_1517448501_2028;
   assign v3_1517448501_2031 = ~v3_1517448501_2032;
   assign v3_1517448501_2032 = ~v3_1517448501_2026 & ~v3_1517448501_2030;
   assign v3_1517448501_2033 = ~v3_1517448501_2034;
   assign v3_1517448501_2034 = ~v3_1517448501_523 & ~v3_1517448501_2028;
   assign v3_1517448501_2035 = v3_1517448501_529 & v3_1517448501_2033;
   assign v3_1517448501_2036 = ~v3_1517448501_2037;
   assign v3_1517448501_2037 = ~v3_1517448501_2031 & ~v3_1517448501_2035;
   assign v3_1517448501_2038 = ~v3_1517448501_2039;
   assign v3_1517448501_2039 = ~v3_1517448501_529 & ~v3_1517448501_2033;
   assign v3_1517448501_2040 = v3_1517448501_532 & v3_1517448501_2038;
   assign v3_1517448501_2041 = ~v3_1517448501_2042;
   assign v3_1517448501_2042 = ~v3_1517448501_2036 & ~v3_1517448501_2040;
   assign v3_1517448501_2043 = v3_1517448501_2021 & ~v3_1517448501_2041;
   assign v3_1517448501_2044 = ~v3_1517448501_2045;
   assign v3_1517448501_2045 = ~v3_1517448501_532 & ~v3_1517448501_2038;
   assign v3_1517448501_2046 = v3_1517448501_2043 & v3_1517448501_2044;
   assign v3_1517448501_2047 = v3_1517448501_557 & v3_1517448501_606;
   assign v3_1517448501_2048 = ~v3_1517448501_2049;
   assign v3_1517448501_2049 = ~v3_1517448501_557 & ~v3_1517448501_606;
   assign v3_1517448501_2050 = v3_1517448501_613 & v3_1517448501_2048;
   assign v3_1517448501_2051 = ~v3_1517448501_2052;
   assign v3_1517448501_2052 = ~v3_1517448501_2047 & ~v3_1517448501_2050;
   assign v3_1517448501_2053 = ~v3_1517448501_2054;
   assign v3_1517448501_2054 = ~v3_1517448501_613 & ~v3_1517448501_2048;
   assign v3_1517448501_2055 = v3_1517448501_623 & v3_1517448501_2053;
   assign v3_1517448501_2056 = ~v3_1517448501_2057;
   assign v3_1517448501_2057 = ~v3_1517448501_2051 & ~v3_1517448501_2055;
   assign v3_1517448501_2058 = ~v3_1517448501_2059;
   assign v3_1517448501_2059 = ~v3_1517448501_623 & ~v3_1517448501_2053;
   assign v3_1517448501_2060 = v3_1517448501_633 & v3_1517448501_2058;
   assign v3_1517448501_2061 = ~v3_1517448501_2062;
   assign v3_1517448501_2062 = ~v3_1517448501_2056 & ~v3_1517448501_2060;
   assign v3_1517448501_2063 = ~v3_1517448501_2064;
   assign v3_1517448501_2064 = ~v3_1517448501_633 & ~v3_1517448501_2058;
   assign v3_1517448501_2065 = v3_1517448501_636 & v3_1517448501_2063;
   assign v3_1517448501_2066 = ~v3_1517448501_2067;
   assign v3_1517448501_2067 = ~v3_1517448501_2061 & ~v3_1517448501_2065;
   assign v3_1517448501_2068 = ~v3_1517448501_2069;
   assign v3_1517448501_2069 = ~v3_1517448501_636 & ~v3_1517448501_2063;
   assign v3_1517448501_2070 = v3_1517448501_641 & v3_1517448501_2068;
   assign v3_1517448501_2071 = ~v3_1517448501_2072;
   assign v3_1517448501_2072 = ~v3_1517448501_2066 & ~v3_1517448501_2070;
   assign v3_1517448501_2073 = v3_1517448501_2046 & ~v3_1517448501_2071;
   assign v3_1517448501_2074 = ~v3_1517448501_2075;
   assign v3_1517448501_2075 = ~v3_1517448501_641 & ~v3_1517448501_2068;
   assign v3_1517448501_2076 = v3_1517448501_2073 & v3_1517448501_2074;
   assign v3_1517448501_2077 = v3_1517448501_666 & v3_1517448501_715;
   assign v3_1517448501_2078 = ~v3_1517448501_2079;
   assign v3_1517448501_2079 = ~v3_1517448501_666 & ~v3_1517448501_715;
   assign v3_1517448501_2080 = v3_1517448501_722 & v3_1517448501_2078;
   assign v3_1517448501_2081 = ~v3_1517448501_2082;
   assign v3_1517448501_2082 = ~v3_1517448501_2077 & ~v3_1517448501_2080;
   assign v3_1517448501_2083 = ~v3_1517448501_2084;
   assign v3_1517448501_2084 = ~v3_1517448501_722 & ~v3_1517448501_2078;
   assign v3_1517448501_2085 = v3_1517448501_732 & v3_1517448501_2083;
   assign v3_1517448501_2086 = ~v3_1517448501_2087;
   assign v3_1517448501_2087 = ~v3_1517448501_2081 & ~v3_1517448501_2085;
   assign v3_1517448501_2088 = ~v3_1517448501_2089;
   assign v3_1517448501_2089 = ~v3_1517448501_732 & ~v3_1517448501_2083;
   assign v3_1517448501_2090 = v3_1517448501_742 & v3_1517448501_2088;
   assign v3_1517448501_2091 = ~v3_1517448501_2092;
   assign v3_1517448501_2092 = ~v3_1517448501_2086 & ~v3_1517448501_2090;
   assign v3_1517448501_2093 = ~v3_1517448501_2094;
   assign v3_1517448501_2094 = ~v3_1517448501_742 & ~v3_1517448501_2088;
   assign v3_1517448501_2095 = v3_1517448501_745 & v3_1517448501_2093;
   assign v3_1517448501_2096 = ~v3_1517448501_2097;
   assign v3_1517448501_2097 = ~v3_1517448501_2091 & ~v3_1517448501_2095;
   assign v3_1517448501_2098 = ~v3_1517448501_2099;
   assign v3_1517448501_2099 = ~v3_1517448501_745 & ~v3_1517448501_2093;
   assign v3_1517448501_2100 = v3_1517448501_750 & v3_1517448501_2098;
   assign v3_1517448501_2101 = ~v3_1517448501_2102;
   assign v3_1517448501_2102 = ~v3_1517448501_2096 & ~v3_1517448501_2100;
   assign v3_1517448501_2103 = v3_1517448501_2076 & ~v3_1517448501_2101;
   assign v3_1517448501_2104 = ~v3_1517448501_2105;
   assign v3_1517448501_2105 = ~v3_1517448501_750 & ~v3_1517448501_2098;
   assign v3_1517448501_2106 = v3_1517448501_2103 & v3_1517448501_2104;
   assign v3_1517448501_2107 = v3_1517448501_798 & v3_1517448501_785;
   assign v3_1517448501_2108 = ~v3_1517448501_2109;
   assign v3_1517448501_2109 = ~v3_1517448501_798 & ~v3_1517448501_785;
   assign v3_1517448501_2110 = v3_1517448501_806 & v3_1517448501_2108;
   assign v3_1517448501_2111 = ~v3_1517448501_2112;
   assign v3_1517448501_2112 = ~v3_1517448501_2107 & ~v3_1517448501_2110;
   assign v3_1517448501_2113 = ~v3_1517448501_2114;
   assign v3_1517448501_2114 = ~v3_1517448501_806 & ~v3_1517448501_2108;
   assign v3_1517448501_2115 = v3_1517448501_815 & v3_1517448501_2113;
   assign v3_1517448501_2116 = ~v3_1517448501_2117;
   assign v3_1517448501_2117 = ~v3_1517448501_2111 & ~v3_1517448501_2115;
   assign v3_1517448501_2118 = ~v3_1517448501_2119;
   assign v3_1517448501_2119 = ~v3_1517448501_815 & ~v3_1517448501_2113;
   assign v3_1517448501_2120 = v3_1517448501_821 & v3_1517448501_2118;
   assign v3_1517448501_2121 = ~v3_1517448501_2122;
   assign v3_1517448501_2122 = ~v3_1517448501_2116 & ~v3_1517448501_2120;
   assign v3_1517448501_2123 = ~v3_1517448501_2124;
   assign v3_1517448501_2124 = ~v3_1517448501_821 & ~v3_1517448501_2118;
   assign v3_1517448501_2125 = v3_1517448501_829 & v3_1517448501_2123;
   assign v3_1517448501_2126 = ~v3_1517448501_2127;
   assign v3_1517448501_2127 = ~v3_1517448501_2121 & ~v3_1517448501_2125;
   assign v3_1517448501_2128 = ~v3_1517448501_2129;
   assign v3_1517448501_2129 = ~v3_1517448501_829 & ~v3_1517448501_2123;
   assign v3_1517448501_2130 = v3_1517448501_836 & v3_1517448501_2128;
   assign v3_1517448501_2131 = ~v3_1517448501_2132;
   assign v3_1517448501_2132 = ~v3_1517448501_2126 & ~v3_1517448501_2130;
   assign v3_1517448501_2133 = ~v3_1517448501_2134;
   assign v3_1517448501_2134 = ~v3_1517448501_836 & ~v3_1517448501_2128;
   assign v3_1517448501_2135 = v3_1517448501_841 & v3_1517448501_2133;
   assign v3_1517448501_2136 = ~v3_1517448501_2137;
   assign v3_1517448501_2137 = ~v3_1517448501_2131 & ~v3_1517448501_2135;
   assign v3_1517448501_2138 = v3_1517448501_2106 & ~v3_1517448501_2136;
   assign v3_1517448501_2139 = ~v3_1517448501_2140;
   assign v3_1517448501_2140 = ~v3_1517448501_841 & ~v3_1517448501_2133;
   assign v3_1517448501_2141 = v3_1517448501_2138 & v3_1517448501_2139;
   assign v3_1517448501_2142 = v3_1517448501_1997 & v3_1517448501_2141;
   assign v3_1517448501_2143 = v3_1517448501_2142 & ~dve_invalid;
   assign v3_1517448501_2144 = 1'b0; 

   // Output Net Assignments
   assign id60 = v3_1517448501_62;

   // Property
   wire prop = !id60;
   wire prop_neg = !prop;
   assert property ( prop );

   // Non-blocking Assignments
   always @ (posedge v3_clock) begin
      v_m_initiator_0 <= v3_1517448501_103;
      v_party_nonce_initiator_0 <= v3_1517448501_134;
      v_m_initiator_1 <= v3_1517448501_145;
      v_party_nonce_initiator_1 <= v3_1517448501_175;
      v_m_responder_0 <= v3_1517448501_267;
      v_party_responder_0 <= v3_1517448501_297;
      v_party_nonce_responder_0 <= v3_1517448501_310;
      v_m_responder_1 <= v3_1517448501_363;
      v_party_responder_1 <= v3_1517448501_393;
      v_party_nonce_responder_1 <= v3_1517448501_406;
      v_kNa <= v3_1517448501_412;
      v_kNb <= v3_1517448501_417;
      v_k_Na_Nb__A <= v3_1517448501_420;
      v_k_Na_A__B <= v3_1517448501_423;
      v_k_Nb__B <= v3_1517448501_428;
      v_m_intruder <= v3_1517448501_441;
      a_start_initiator_0 <= ~v3_1517448501_445;
      a_wait_resp_initiator_0 <= v3_1517448501_457;
      a_got_resp_initiator_0 <= v3_1517448501_470;
      a_commited_initiator_0 <= v3_1517448501_477;
      a_finished_initiator_0 <= v3_1517448501_483;
      a_corrupted_initiator_0 <= v3_1517448501_486;
      a_start_initiator_1 <= ~v3_1517448501_491;
      a_wait_resp_initiator_1 <= v3_1517448501_503;
      a_got_resp_initiator_1 <= v3_1517448501_516;
      a_commited_initiator_1 <= v3_1517448501_523;
      a_finished_initiator_1 <= v3_1517448501_529;
      a_corrupted_initiator_1 <= v3_1517448501_532;
      a_start_responder_0 <= ~v3_1517448501_557;
      a_got_msg_responder_0 <= v3_1517448501_606;
      a_send_reply_responder_0 <= v3_1517448501_613;
      a_wait_resp_responder_0 <= v3_1517448501_623;
      a_got_resp_responder_0 <= v3_1517448501_633;
      a_finished_responder_0 <= v3_1517448501_636;
      a_corrupted_responder_0 <= v3_1517448501_641;
      a_start_responder_1 <= ~v3_1517448501_666;
      a_got_msg_responder_1 <= v3_1517448501_715;
      a_send_reply_responder_1 <= v3_1517448501_722;
      a_wait_resp_responder_1 <= v3_1517448501_732;
      a_got_resp_responder_1 <= v3_1517448501_742;
      a_finished_responder_1 <= v3_1517448501_745;
      a_corrupted_responder_1 <= v3_1517448501_750;
      a_q <= ~v3_1517448501_785;
      a_got3 <= v3_1517448501_798;
      a_c1 <= v3_1517448501_806;
      a_c2 <= v3_1517448501_815;
      a_d1 <= v3_1517448501_821;
      a_got2 <= v3_1517448501_829;
      a_e1 <= v3_1517448501_836;
      a_f1 <= v3_1517448501_841;
      dve_invalid <= ~v3_1517448501_2143;
   end
endmodule
